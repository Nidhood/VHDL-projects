LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE texturas IS

	TYPE ImageMatrix IS ARRAY (NATURAL RANGE <>, NATURAL RANGE <>) OF STD_logic_vector(7 DOWNTO 0);

	-------------------------------------------------------------------------------------------
	------------------------------- Moto Derecha ----------------------------------------------
	-------------------------------------------------------------------------------------------

CONSTANT MotoPlantilla_DerechaR : ImageMatrix(0 TO 49, 0 TO 49) := (
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"7F" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"0C" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"7F" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"7F" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"7F" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"7F" , x"00" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"00" , x"7F" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"00" , x"7F" , x"FF" , x"FF" ),
( x"FF" , x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"FF" ),
( x"FF" , x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"FF" ),
( x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" ),
( x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" ),
( x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" ),
( x"FF" , x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"FF" ),
( x"FF" , x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"FF" ),
( x"FF" , x"FF" , x"7F" , x"00" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"00" , x"7F" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"00" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"00" , x"7F" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"7F" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"7F" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"7F" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"7F" , x"7F" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"7F" , x"7F" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ) 
);

CONSTANT MotoPlantilla_DerechaG : ImageMatrix(0 TO 49, 0 TO 49) := (
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"7F" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"C7" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"7F" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"7F" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"7F" , x"00" , x"00" ),
( x"00" , x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"00" ),
( x"00" , x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"00" ),
( x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" ),
( x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" ),
( x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" ),
( x"00" , x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"00" ),
( x"00" , x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"00" ),
( x"00" , x"00" , x"7F" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"7F" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ) 
);

CONSTANT MotoPlantilla_DerechaB : ImageMatrix(0 TO 49, 0 TO 49) := (
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"7F" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"FA" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"7F" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"7F" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"7F" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"7F" , x"00" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"00" , x"7F" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"00" , x"7F" , x"DC" , x"DC" ),
( x"DC" , x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"DC" ),
( x"DC" , x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"DC" ),
( x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" ),
( x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" ),
( x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" ),
( x"DC" , x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"DC" ),
( x"DC" , x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"DC" ),
( x"DC" , x"DC" , x"7F" , x"00" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"00" , x"7F" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"00" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"00" , x"7F" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"7F" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"7F" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"7F" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"7F" , x"7F" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"7F" , x"7F" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ) 
);



	-------------------------------------------------------------------------------------------
	------------------------------------ Vidas ------------------------------------------
	-------------------------------------------------------------------------------------------	
	
CONSTANT VidasR : ImageMatrix(0 TO 49, 0 TO 34) := (
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"0C" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"0C" , x"FF" , x"FF" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"0C" , x"FF" , x"FF" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"0C" , x"FF" , x"FF" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"0C" , x"FF" , x"FF" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"FF" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"00" , x"FF" , x"00" , x"00" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"00" , x"FF" , x"00" , x"00" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"0C" , x"0C" , x"00" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"0C" , x"00" , x"00" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"00" , x"00" , x"0C" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"0C" , x"0C" , x"0C" , x"0C" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"0C" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ) 
);

CONSTANT VidasG : ImageMatrix(0 TO 49, 0 TO 34) := (
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"C7" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"C7" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"C7" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"C7" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"C7" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"C7" , x"C7" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"C7" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ),
( x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" ) 
);

CONSTANT VidasB : ImageMatrix(0 TO 49, 0 TO 34) := (
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"7F" , x"7F" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"FA" , x"DC" , x"DC" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"FA" , x"DC" , x"DC" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"FA" , x"DC" , x"DC" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"FA" , x"DC" , x"DC" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"7F" , x"7F" , x"00" , x"DC" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"00" , x"DC" , x"00" , x"00" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"00" , x"DC" , x"00" , x"00" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"FA" , x"FA" , x"00" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"FA" , x"00" , x"00" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"00" , x"00" , x"FA" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"FA" , x"FA" , x"FA" , x"FA" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"FA" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"00" , x"00" , x"00" , x"00" , x"00" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ),
( x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" , x"DC" ) 
);

---------------------------------------------------------------

END PACKAGE texturas;

-------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------------

PACKAGE BODY texturas IS

END texturas;