---------------------------------------------------------------------------------
--                                                                             -- 
--    Two shifter: Shifts the input one times to the left, to multiply by 2.   --
--    Author: Ivan Dario Orozco Ibanez                                         --
--                                                                             --
---------------------------------------------------------------------------------