LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY fpga03 IS
    PORT (
        bin : IN STD_LOGIC_VECTOR(10 DOWNTO 0);
        led : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
    );
END ENTITY fpga03;

ARCHITECTURE functional OF fpga03 IS
BEGIN

    WITH bin SELECT
        led <=
        "0000000001" WHEN "10000000001",
        "0000000010" WHEN "00000000010",
        "0000000100" WHEN "10000000100",
        "0000001000" WHEN "00000001000",
        "0000010000" WHEN "10000010000",
        "0000100000" WHEN "00000100000",
        "0001000000" WHEN "10001000000",
        "0010000000" WHEN "00010000000",
        "0100000000" WHEN "10100000000",
        "1000000000" WHEN "01000000000",
        "0000000000" WHEN OTHERS;

END ARCHITECTURE functional;