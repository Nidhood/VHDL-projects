LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

PACKAGE texturas IS

	TYPE ImageMatrix IS ARRAY (NATURAL RANGE <>, NATURAL RANGE <>) OF STD_logic_vector(7 DOWNTO 0);

	-------------------------------------------------------------------------------------------
	------------------------------- Moto Derecha ----------------------------------------------
	-------------------------------------------------------------------------------------------

CONSTANT MotoPlantilla_DerechaR : ImageMatrix(0 TO 39, 0 TO 39) := (
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"32" , x"32" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"32" , x"32" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"E1" , x"E1" , x"00" , x"00" , x"00" , x"32" , x"32" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"32" , x"32" , x"32" , x"32" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"00" , x"32" , x"32" , x"32" , x"00" , x"32" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"00" , x"32" , x"32" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"00" , x"00" , x"00" , x"32" , x"32" , x"32" , x"32" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"32" , x"32" , x"32" , x"00" , x"54" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"80" , x"00" , x"00" , x"E1" , x"E1" , x"00" , x"00" , x"00" , x"00" , x"00" , x"32" , x"32" , x"00" , x"00" , x"00" , x"32" , x"32" , x"32" , x"00" , x"00" , x"54" , x"54" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"00" , x"00" , x"E1" , x"E1" ),
( x"E1" , x"00" , x"80" , x"80" , x"80" , x"00" , x"00" , x"00" , x"80" , x"80" , x"80" , x"00" , x"E1" , x"00" , x"54" , x"54" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"32" , x"32" , x"32" , x"00" , x"54" , x"54" , x"54" , x"54" , x"00" , x"00" , x"00" , x"00" , x"80" , x"80" , x"80" , x"00" , x"E1" ),
( x"E1" , x"00" , x"80" , x"80" , x"00" , x"00" , x"00" , x"00" , x"00" , x"80" , x"80" , x"00" , x"00" , x"54" , x"54" , x"00" , x"00" , x"00" , x"00" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"E1" , x"00" , x"00" , x"54" , x"54" , x"54" , x"E1" , x"00" , x"00" , x"00" , x"80" , x"80" , x"00" , x"E1" ),
( x"00" , x"80" , x"80" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"80" , x"00" , x"00" , x"54" , x"00" , x"54" , x"54" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"E1" , x"00" , x"00" , x"00" , x"54" , x"54" , x"54" , x"E1" , x"E1" , x"00" , x"00" , x"80" , x"80" , x"00" ),
( x"00" , x"80" , x"00" , x"00" , x"E1" , x"E1" , x"00" , x"00" , x"54" , x"54" , x"54" , x"54" , x"54" , x"00" , x"54" , x"54" , x"00" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"E1" , x"00" , x"80" , x"00" , x"54" , x"54" , x"54" , x"00" , x"00" , x"E1" , x"00" , x"00" , x"80" , x"00" ),
( x"00" , x"80" , x"00" , x"00" , x"E1" , x"00" , x"E1" , x"00" , x"54" , x"54" , x"54" , x"54" , x"54" , x"00" , x"54" , x"00" , x"00" , x"00" , x"32" , x"32" , x"32" , x"00" , x"32" , x"32" , x"32" , x"00" , x"E1" , x"00" , x"80" , x"00" , x"00" , x"E1" , x"00" , x"E1" , x"00" , x"E1" , x"00" , x"00" , x"80" , x"00" ),
( x"00" , x"80" , x"00" , x"00" , x"E1" , x"00" , x"00" , x"00" , x"54" , x"54" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"E1" , x"00" , x"80" , x"00" , x"00" , x"E1" , x"00" , x"00" , x"00" , x"E1" , x"00" , x"00" , x"80" , x"00" ),
( x"00" , x"80" , x"80" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"80" , x"80" , x"00" , x"00" , x"32" , x"32" , x"32" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"E1" , x"00" , x"80" , x"80" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"80" , x"80" , x"00" ),
( x"E1" , x"00" , x"80" , x"80" , x"00" , x"00" , x"00" , x"00" , x"00" , x"80" , x"80" , x"00" , x"E1" , x"00" , x"00" , x"00" , x"00" , x"32" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"E1" , x"E1" , x"00" , x"80" , x"80" , x"00" , x"00" , x"00" , x"00" , x"00" , x"80" , x"80" , x"00" , x"E1" ),
( x"E1" , x"00" , x"80" , x"80" , x"80" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"32" , x"00" , x"E1" , x"E1" , x"00" , x"80" , x"80" , x"80" , x"00" , x"00" , x"00" , x"80" , x"80" , x"80" , x"00" , x"E1" ),
( x"E1" , x"E1" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"80" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"80" , x"00" , x"00" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"00" , x"00" , x"00" , x"00" , x"00" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ),
( x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" , x"E1" ) 
);

CONSTANT MotoPlantilla_DerechaG : ImageMatrix(0 TO 39, 0 TO 39) := (
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"00" , x"00" , x"00" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"82" , x"82" , x"00" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"07" , x"07" , x"07" , x"07" , x"00" , x"82" , x"82" , x"00" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"00" , x"00" , x"00" , x"00" , x"00" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"07" , x"07" , x"00" , x"00" , x"00" , x"82" , x"82" , x"00" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"00" , x"82" , x"82" , x"82" , x"82" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"00" , x"82" , x"82" , x"82" , x"00" , x"82" , x"00" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"00" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"00" , x"82" , x"82" , x"00" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"00" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"00" , x"00" , x"00" , x"82" , x"82" , x"82" , x"82" , x"00" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"00" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"00" , x"00" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"00" , x"00" , x"00" , x"00" , x"00" , x"07" , x"07" , x"07" , x"07" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"82" , x"82" , x"82" , x"00" , x"54" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"80" , x"00" , x"00" , x"07" , x"07" , x"00" , x"00" , x"00" , x"00" , x"00" , x"82" , x"82" , x"00" , x"00" , x"00" , x"82" , x"82" , x"82" , x"00" , x"00" , x"54" , x"54" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"00" , x"00" , x"07" , x"07" ),
( x"07" , x"00" , x"80" , x"80" , x"80" , x"00" , x"00" , x"00" , x"80" , x"80" , x"80" , x"00" , x"07" , x"00" , x"54" , x"54" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"82" , x"82" , x"82" , x"00" , x"54" , x"54" , x"54" , x"54" , x"00" , x"00" , x"00" , x"00" , x"80" , x"80" , x"80" , x"00" , x"07" ),
( x"07" , x"00" , x"80" , x"80" , x"00" , x"00" , x"00" , x"00" , x"00" , x"80" , x"80" , x"00" , x"00" , x"54" , x"54" , x"00" , x"00" , x"00" , x"00" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"07" , x"00" , x"00" , x"54" , x"54" , x"54" , x"07" , x"00" , x"00" , x"00" , x"80" , x"80" , x"00" , x"07" ),
( x"00" , x"80" , x"80" , x"00" , x"00" , x"07" , x"07" , x"07" , x"00" , x"00" , x"80" , x"00" , x"00" , x"54" , x"00" , x"54" , x"54" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"07" , x"00" , x"00" , x"00" , x"54" , x"54" , x"54" , x"07" , x"07" , x"00" , x"00" , x"80" , x"80" , x"00" ),
( x"00" , x"80" , x"00" , x"00" , x"07" , x"07" , x"00" , x"00" , x"54" , x"54" , x"54" , x"54" , x"54" , x"00" , x"54" , x"54" , x"00" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"07" , x"00" , x"80" , x"00" , x"54" , x"54" , x"54" , x"00" , x"00" , x"07" , x"00" , x"00" , x"80" , x"00" ),
( x"00" , x"80" , x"00" , x"00" , x"07" , x"00" , x"07" , x"00" , x"54" , x"54" , x"54" , x"54" , x"54" , x"00" , x"54" , x"00" , x"00" , x"00" , x"82" , x"82" , x"82" , x"00" , x"82" , x"82" , x"82" , x"00" , x"07" , x"00" , x"80" , x"00" , x"00" , x"07" , x"00" , x"07" , x"00" , x"07" , x"00" , x"00" , x"80" , x"00" ),
( x"00" , x"80" , x"00" , x"00" , x"07" , x"00" , x"00" , x"00" , x"54" , x"54" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"07" , x"00" , x"80" , x"00" , x"00" , x"07" , x"00" , x"00" , x"00" , x"07" , x"00" , x"00" , x"80" , x"00" ),
( x"00" , x"80" , x"80" , x"00" , x"00" , x"07" , x"07" , x"07" , x"00" , x"00" , x"80" , x"80" , x"00" , x"00" , x"82" , x"82" , x"82" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"07" , x"00" , x"80" , x"80" , x"00" , x"00" , x"07" , x"07" , x"07" , x"00" , x"00" , x"80" , x"80" , x"00" ),
( x"07" , x"00" , x"80" , x"80" , x"00" , x"00" , x"00" , x"00" , x"00" , x"80" , x"80" , x"00" , x"07" , x"00" , x"00" , x"00" , x"00" , x"82" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"07" , x"07" , x"00" , x"80" , x"80" , x"00" , x"00" , x"00" , x"00" , x"00" , x"80" , x"80" , x"00" , x"07" ),
( x"07" , x"00" , x"80" , x"80" , x"80" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"00" , x"07" , x"07" , x"07" , x"07" , x"07" , x"00" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"82" , x"00" , x"07" , x"07" , x"00" , x"80" , x"80" , x"80" , x"00" , x"00" , x"00" , x"80" , x"80" , x"80" , x"00" , x"07" ),
( x"07" , x"07" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"80" , x"00" , x"00" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"07" , x"07" , x"07" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"80" , x"00" , x"00" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"00" , x"00" , x"00" , x"00" , x"00" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"00" , x"00" , x"00" , x"00" , x"00" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ),
( x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" , x"07" ) 
);

CONSTANT MotoPlantilla_DerechaB : ImageMatrix(0 TO 39, 0 TO 39) := (
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"F6" , x"F6" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"F6" , x"F6" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"F6" , x"F6" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"00" , x"F6" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"00" , x"F6" , x"F6" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"00" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"F6" , x"F6" , x"F6" , x"00" , x"54" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"80" , x"00" , x"00" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"F6" , x"F6" , x"00" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"00" , x"00" , x"54" , x"54" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"00" , x"00" , x"FF" , x"FF" ),
( x"FF" , x"00" , x"80" , x"80" , x"80" , x"00" , x"00" , x"00" , x"80" , x"80" , x"80" , x"00" , x"FF" , x"00" , x"54" , x"54" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"00" , x"54" , x"54" , x"54" , x"54" , x"00" , x"00" , x"00" , x"00" , x"80" , x"80" , x"80" , x"00" , x"FF" ),
( x"FF" , x"00" , x"80" , x"80" , x"00" , x"00" , x"00" , x"00" , x"00" , x"80" , x"80" , x"00" , x"00" , x"54" , x"54" , x"00" , x"00" , x"00" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"FF" , x"00" , x"00" , x"54" , x"54" , x"54" , x"FF" , x"00" , x"00" , x"00" , x"80" , x"80" , x"00" , x"FF" ),
( x"00" , x"80" , x"80" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"80" , x"00" , x"00" , x"54" , x"00" , x"54" , x"54" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"FF" , x"00" , x"00" , x"00" , x"54" , x"54" , x"54" , x"FF" , x"FF" , x"00" , x"00" , x"80" , x"80" , x"00" ),
( x"00" , x"80" , x"00" , x"00" , x"FF" , x"FF" , x"00" , x"00" , x"54" , x"54" , x"54" , x"54" , x"54" , x"00" , x"54" , x"54" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"FF" , x"00" , x"80" , x"00" , x"54" , x"54" , x"54" , x"00" , x"00" , x"FF" , x"00" , x"00" , x"80" , x"00" ),
( x"00" , x"80" , x"00" , x"00" , x"FF" , x"00" , x"FF" , x"00" , x"54" , x"54" , x"54" , x"54" , x"54" , x"00" , x"54" , x"00" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"00" , x"F6" , x"F6" , x"F6" , x"00" , x"FF" , x"00" , x"80" , x"00" , x"00" , x"FF" , x"00" , x"FF" , x"00" , x"FF" , x"00" , x"00" , x"80" , x"00" ),
( x"00" , x"80" , x"00" , x"00" , x"FF" , x"00" , x"00" , x"00" , x"54" , x"54" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"FF" , x"00" , x"80" , x"00" , x"00" , x"FF" , x"00" , x"00" , x"00" , x"FF" , x"00" , x"00" , x"80" , x"00" ),
( x"00" , x"80" , x"80" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"80" , x"80" , x"00" , x"00" , x"F6" , x"F6" , x"F6" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"FF" , x"00" , x"80" , x"80" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"80" , x"80" , x"00" ),
( x"FF" , x"00" , x"80" , x"80" , x"00" , x"00" , x"00" , x"00" , x"00" , x"80" , x"80" , x"00" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"F6" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"FF" , x"FF" , x"00" , x"80" , x"80" , x"00" , x"00" , x"00" , x"00" , x"00" , x"80" , x"80" , x"00" , x"FF" ),
( x"FF" , x"00" , x"80" , x"80" , x"80" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"00" , x"FF" , x"FF" , x"00" , x"80" , x"80" , x"80" , x"00" , x"00" , x"00" , x"80" , x"80" , x"80" , x"00" , x"FF" ),
( x"FF" , x"FF" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"80" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"80" , x"80" , x"80" , x"80" , x"80" , x"00" , x"00" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"00" , x"00" , x"00" , x"00" , x"00" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ) 
);


	-------------------------------------------------------------------------------------------
	------------------------------------ Titulo Tron ------------------------------------------
	-------------------------------------------------------------------------------------------	
	
	
	CONSTANT Plantilla_TronR : ImageMatrix(0 TO 99, 0 TO 99) := (
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"FD" , x"FE" , x"FF" , x"FF" , x"FE" , x"FD" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FC" , x"FD" , x"FE" , x"FD" , x"FD" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FD" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FC" , x"FF" , x"FF" , x"FF" , x"FD" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FD" , x"FB" , x"FB" , x"FD" , x"FD" , x"FE" , x"FD" , x"FD" , x"FE" , x"FD" , x"FE" , x"FE" , x"FE" , x"FD" , x"FB" , x"F9" , x"F8" , x"FB" , x"FD" , x"FA" , x"FA" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"F9" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"A2" , x"63" , x"5D" , x"5F" , x"64" , x"68" , x"71" , x"94" , x"F0" , x"FF" , x"FF" , x"FA" , x"AC" , x"78" , x"61" , x"5B" , x"5B" , x"58" , x"59" , x"5B" , x"5D" , x"5E" , x"5D" , x"5D" , x"5E" , x"5B" , x"5B" , x"5E" , x"5E" , x"5B" , x"5A" , x"56" , x"55" , x"5A" , x"5B" , x"56" , x"56" , x"62" , x"84" , x"C1" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FE" , x"BD" , x"84" , x"69" , x"71" , x"A4" , x"EE" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"DC" , x"7F" , x"60" , x"A1" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"F7" , x"8E" , x"5E" , x"55" , x"61" , x"7D" , x"E4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FD" , x"FF" , x"B8" , x"34" , x"37" , x"37" , x"36" , x"36" , x"36" , x"36" , x"39" , x"7F" , x"FF" , x"F8" , x"6E" , x"35" , x"37" , x"36" , x"36" , x"36" , x"36" , x"36" , x"35" , x"35" , x"35" , x"35" , x"35" , x"36" , x"36" , x"36" , x"35" , x"35" , x"35" , x"35" , x"35" , x"35" , x"35" , x"36" , x"36" , x"35" , x"36" , x"36" , x"34" , x"81" , x"FA" , x"FD" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"EC" , x"6D" , x"31" , x"35" , x"37" , x"35" , x"34" , x"51" , x"CF" , x"FF" , x"FD" , x"FF" , x"FF" , x"FE" , x"FE" , x"FA" , x"57" , x"38" , x"37" , x"37" , x"C5" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"A3" , x"36" , x"37" , x"36" , x"37" , x"39" , x"65" , x"FD" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FD" , x"FF" , x"73" , x"57" , x"77" , x"6F" , x"72" , x"72" , x"72" , x"75" , x"6B" , x"3F" , x"F8" , x"A4" , x"37" , x"5C" , x"71" , x"72" , x"71" , x"71" , x"71" , x"70" , x"6F" , x"6F" , x"71" , x"6F" , x"6F" , x"72" , x"71" , x"70" , x"71" , x"71" , x"6F" , x"6F" , x"6F" , x"6F" , x"6F" , x"70" , x"71" , x"70" , x"72" , x"6D" , x"4C" , x"36" , x"83" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"F3" , x"59" , x"36" , x"4A" , x"69" , x"71" , x"6D" , x"56" , x"39" , x"3E" , x"D1" , x"FF" , x"FD" , x"FF" , x"FC" , x"FF" , x"CF" , x"40" , x"6E" , x"79" , x"61" , x"75" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"65" , x"59" , x"75" , x"6E" , x"72" , x"6B" , x"39" , x"DC" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"5D" , x"84" , x"99" , x"93" , x"95" , x"95" , x"95" , x"95" , x"97" , x"4E" , x"CB" , x"58" , x"5F" , x"94" , x"92" , x"95" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"95" , x"95" , x"96" , x"8E" , x"5E" , x"30" , x"C6" , x"FF" , x"FC" , x"FF" , x"FF" , x"FD" , x"FF" , x"7A" , x"38" , x"62" , x"8B" , x"94" , x"93" , x"94" , x"91" , x"73" , x"3F" , x"4A" , x"F0" , x"FD" , x"FE" , x"FC" , x"FF" , x"A7" , x"67" , x"9D" , x"96" , x"86" , x"4B" , x"F6" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FE" , x"55" , x"85" , x"99" , x"94" , x"93" , x"97" , x"56" , x"B5" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"FB" , x"57" , x"89" , x"83" , x"82" , x"84" , x"83" , x"83" , x"80" , x"8D" , x"5D" , x"6C" , x"4C" , x"8B" , x"8E" , x"7F" , x"82" , x"82" , x"83" , x"82" , x"83" , x"83" , x"83" , x"83" , x"83" , x"83" , x"83" , x"82" , x"83" , x"83" , x"83" , x"83" , x"83" , x"83" , x"83" , x"83" , x"83" , x"82" , x"83" , x"84" , x"86" , x"93" , x"92" , x"51" , x"64" , x"FF" , x"FE" , x"FF" , x"FC" , x"FF" , x"C1" , x"33" , x"65" , x"93" , x"92" , x"89" , x"83" , x"85" , x"8E" , x"95" , x"79" , x"3D" , x"87" , x"FF" , x"FD" , x"FC" , x"FF" , x"92" , x"7B" , x"8E" , x"81" , x"8E" , x"4C" , x"CA" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F7" , x"57" , x"8C" , x"84" , x"85" , x"7F" , x"8F" , x"6E" , x"A3" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F6" , x"56" , x"82" , x"41" , x"3E" , x"3D" , x"3D" , x"41" , x"39" , x"6C" , x"66" , x"23" , x"62" , x"94" , x"56" , x"3E" , x"3F" , x"40" , x"40" , x"3F" , x"40" , x"41" , x"41" , x"41" , x"41" , x"41" , x"41" , x"41" , x"40" , x"40" , x"41" , x"40" , x"3F" , x"40" , x"3E" , x"3E" , x"3F" , x"40" , x"3F" , x"3E" , x"42" , x"63" , x"92" , x"80" , x"39" , x"DB" , x"FF" , x"FC" , x"FE" , x"F8" , x"4B" , x"56" , x"93" , x"8C" , x"65" , x"46" , x"41" , x"43" , x"5A" , x"84" , x"98" , x"6C" , x"38" , x"DE" , x"FE" , x"FA" , x"FF" , x"82" , x"80" , x"52" , x"37" , x"7F" , x"6E" , x"91" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F4" , x"61" , x"7F" , x"3C" , x"40" , x"39" , x"5F" , x"75" , x"9E" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F5" , x"53" , x"84" , x"3D" , x"32" , x"33" , x"3A" , x"52" , x"40" , x"6D" , x"68" , x"30" , x"81" , x"71" , x"31" , x"33" , x"30" , x"2F" , x"2F" , x"30" , x"2F" , x"30" , x"30" , x"30" , x"30" , x"2F" , x"2F" , x"2F" , x"2F" , x"30" , x"30" , x"30" , x"2F" , x"2F" , x"2F" , x"2F" , x"2F" , x"2F" , x"30" , x"30" , x"33" , x"33" , x"60" , x"99" , x"57" , x"97" , x"FF" , x"F9" , x"FF" , x"AC" , x"3D" , x"84" , x"8D" , x"52" , x"33" , x"32" , x"31" , x"32" , x"34" , x"42" , x"80" , x"92" , x"4F" , x"7D" , x"FF" , x"FB" , x"FF" , x"74" , x"84" , x"54" , x"43" , x"64" , x"85" , x"5F" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F2" , x"60" , x"7E" , x"3B" , x"5C" , x"3F" , x"5A" , x"78" , x"9D" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F4" , x"53" , x"86" , x"5A" , x"D0" , x"D5" , x"DD" , x"F4" , x"AB" , x"6E" , x"68" , x"41" , x"8D" , x"4C" , x"79" , x"BD" , x"C7" , x"C1" , x"BE" , x"BB" , x"BA" , x"B5" , x"AB" , x"A9" , x"AF" , x"B6" , x"B9" , x"B8" , x"B6" , x"B1" , x"AC" , x"B0" , x"BA" , x"C4" , x"CA" , x"C9" , x"C5" , x"C3" , x"BF" , x"B8" , x"B2" , x"6B" , x"38" , x"83" , x"7C" , x"60" , x"FF" , x"FE" , x"F9" , x"4B" , x"68" , x"98" , x"5B" , x"33" , x"67" , x"A3" , x"AD" , x"A3" , x"75" , x"2F" , x"46" , x"8F" , x"7B" , x"3C" , x"E6" , x"FF" , x"FF" , x"6B" , x"85" , x"66" , x"C6" , x"4F" , x"8E" , x"4A" , x"DC" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F0" , x"61" , x"81" , x"6A" , x"FA" , x"AC" , x"5B" , x"79" , x"9D" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F3" , x"55" , x"85" , x"76" , x"FF" , x"FF" , x"FF" , x"FF" , x"C7" , x"6D" , x"65" , x"54" , x"85" , x"55" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"67" , x"58" , x"8D" , x"43" , x"E6" , x"FF" , x"B7" , x"3A" , x"8B" , x"7A" , x"36" , x"90" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"B7" , x"31" , x"5E" , x"99" , x"53" , x"98" , x"FF" , x"FF" , x"65" , x"84" , x"63" , x"FF" , x"61" , x"84" , x"66" , x"9C" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F0" , x"60" , x"81" , x"80" , x"FF" , x"CF" , x"57" , x"78" , x"9F" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F3" , x"55" , x"86" , x"76" , x"FC" , x"FB" , x"FB" , x"FE" , x"C0" , x"6D" , x"63" , x"65" , x"76" , x"8D" , x"FF" , x"F9" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FA" , x"FF" , x"D8" , x"3C" , x"89" , x"52" , x"BC" , x"FF" , x"65" , x"5E" , x"95" , x"49" , x"6A" , x"FF" , x"FC" , x"FA" , x"FD" , x"FB" , x"FA" , x"FF" , x"99" , x"39" , x"87" , x"79" , x"54" , x"FC" , x"FF" , x"60" , x"84" , x"5D" , x"FE" , x"8F" , x"6B" , x"80" , x"5C" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F0" , x"62" , x"81" , x"7F" , x"FE" , x"CE" , x"58" , x"79" , x"9F" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F3" , x"56" , x"86" , x"78" , x"FD" , x"FB" , x"FA" , x"FC" , x"C2" , x"6D" , x"62" , x"71" , x"63" , x"B6" , x"FE" , x"FD" , x"FD" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FD" , x"FD" , x"FD" , x"FD" , x"FC" , x"FD" , x"FD" , x"FD" , x"FD" , x"FE" , x"FE" , x"FE" , x"FD" , x"FE" , x"FE" , x"FF" , x"FE" , x"FE" , x"FE" , x"FC" , x"FD" , x"69" , x"78" , x"6A" , x"9B" , x"F6" , x"38" , x"80" , x"78" , x"3E" , x"E5" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FB" , x"FB" , x"4E" , x"5A" , x"91" , x"42" , x"D0" , x"FF" , x"59" , x"84" , x"5A" , x"FF" , x"C8" , x"4B" , x"8E" , x"45" , x"D8" , x"FF" , x"FD" , x"FF" , x"FF" , x"FE" , x"FF" , x"F1" , x"62" , x"81" , x"7F" , x"FF" , x"CF" , x"58" , x"79" , x"A0" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F3" , x"56" , x"86" , x"72" , x"FF" , x"FF" , x"FF" , x"FF" , x"CB" , x"6C" , x"64" , x"75" , x"55" , x"D5" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"AE" , x"66" , x"78" , x"88" , x"C3" , x"44" , x"93" , x"52" , x"94" , x"FF" , x"FF" , x"DC" , x"7E" , x"5E" , x"7A" , x"DA" , x"FF" , x"FF" , x"BC" , x"39" , x"8B" , x"60" , x"8D" , x"FF" , x"57" , x"83" , x"5D" , x"F9" , x"F6" , x"49" , x"87" , x"5F" , x"99" , x"FF" , x"FC" , x"FF" , x"FF" , x"FE" , x"FF" , x"F2" , x"61" , x"81" , x"7F" , x"FF" , x"D0" , x"58" , x"79" , x"A1" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F3" , x"53" , x"84" , x"46" , x"78" , x"81" , x"88" , x"9A" , x"6D" , x"6E" , x"66" , x"79" , x"52" , x"E4" , x"FF" , x"FF" , x"E1" , x"97" , x"88" , x"7F" , x"7E" , x"80" , x"7C" , x"73" , x"72" , x"7C" , x"84" , x"80" , x"77" , x"74" , x"6F" , x"6D" , x"6D" , x"71" , x"73" , x"72" , x"66" , x"5F" , x"67" , x"6A" , x"6B" , x"76" , x"98" , x"72" , x"5A" , x"80" , x"80" , x"8E" , x"63" , x"88" , x"3F" , x"E7" , x"FF" , x"CC" , x"3D" , x"36" , x"35" , x"36" , x"3E" , x"CD" , x"FF" , x"FD" , x"56" , x"6F" , x"7D" , x"5A" , x"FF" , x"5B" , x"83" , x"5F" , x"F2" , x"FF" , x"79" , x"70" , x"7A" , x"5B" , x"FF" , x"FD" , x"FF" , x"FF" , x"FE" , x"FF" , x"F2" , x"61" , x"81" , x"7B" , x"FF" , x"CF" , x"58" , x"79" , x"A1" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F4" , x"54" , x"82" , x"3A" , x"34" , x"36" , x"35" , x"36" , x"30" , x"69" , x"6A" , x"79" , x"51" , x"EA" , x"FF" , x"F6" , x"53" , x"34" , x"34" , x"34" , x"35" , x"36" , x"35" , x"34" , x"34" , x"34" , x"35" , x"35" , x"35" , x"34" , x"34" , x"34" , x"34" , x"34" , x"35" , x"35" , x"35" , x"35" , x"34" , x"34" , x"35" , x"35" , x"35" , x"34" , x"4C" , x"81" , x"59" , x"51" , x"7D" , x"6E" , x"74" , x"FF" , x"E5" , x"40" , x"38" , x"58" , x"66" , x"5A" , x"3D" , x"46" , x"EB" , x"FE" , x"AB" , x"50" , x"8C" , x"47" , x"EC" , x"64" , x"84" , x"60" , x"F3" , x"FF" , x"BC" , x"52" , x"8D" , x"40" , x"DE" , x"FF" , x"FD" , x"FF" , x"FE" , x"FF" , x"F2" , x"61" , x"81" , x"79" , x"FF" , x"CE" , x"58" , x"79" , x"A2" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F6" , x"52" , x"85" , x"5D" , x"5C" , x"5D" , x"5C" , x"5D" , x"54" , x"77" , x"69" , x"7A" , x"51" , x"EA" , x"FF" , x"B7" , x"38" , x"5A" , x"5C" , x"5B" , x"5C" , x"5C" , x"5B" , x"5A" , x"59" , x"59" , x"59" , x"5A" , x"59" , x"5A" , x"5B" , x"5C" , x"5A" , x"58" , x"5A" , x"5A" , x"5A" , x"5A" , x"59" , x"59" , x"59" , x"5A" , x"5B" , x"57" , x"61" , x"80" , x"2A" , x"34" , x"89" , x"4F" , x"BF" , x"FF" , x"76" , x"37" , x"6E" , x"91" , x"93" , x"93" , x"79" , x"3C" , x"82" , x"FF" , x"ED" , x"46" , x"8B" , x"53" , x"C3" , x"6C" , x"84" , x"5F" , x"F6" , x"FF" , x"F2" , x"4B" , x"8B" , x"59" , x"A0" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"F2" , x"62" , x"81" , x"77" , x"FF" , x"CF" , x"58" , x"79" , x"A3" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"FC" , x"56" , x"89" , x"91" , x"8E" , x"8F" , x"8F" , x"8E" , x"8F" , x"95" , x"60" , x"7D" , x"51" , x"ED" , x"FF" , x"76" , x"60" , x"98" , x"8F" , x"8E" , x"8F" , x"8E" , x"90" , x"92" , x"92" , x"92" , x"92" , x"91" , x"91" , x"92" , x"90" , x"8E" , x"91" , x"92" , x"90" , x"90" , x"90" , x"90" , x"90" , x"90" , x"90" , x"90" , x"90" , x"91" , x"93" , x"81" , x"2D" , x"4C" , x"8A" , x"50" , x"FA" , x"EA" , x"33" , x"63" , x"97" , x"8F" , x"87" , x"8E" , x"97" , x"6C" , x"39" , x"E6" , x"FF" , x"72" , x"79" , x"6C" , x"9D" , x"73" , x"84" , x"60" , x"F7" , x"FF" , x"FF" , x"77" , x"76" , x"76" , x"65" , x"FF" , x"FE" , x"FF" , x"FE" , x"FF" , x"F2" , x"61" , x"81" , x"79" , x"FF" , x"CF" , x"58" , x"79" , x"A3" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FE" , x"FF" , x"62" , x"76" , x"95" , x"8E" , x"90" , x"90" , x"90" , x"92" , x"88" , x"4C" , x"80" , x"52" , x"F2" , x"FF" , x"54" , x"7F" , x"93" , x"8C" , x"8F" , x"8F" , x"90" , x"8F" , x"8E" , x"8F" , x"8F" , x"8F" , x"8F" , x"8E" , x"8E" , x"8F" , x"90" , x"90" , x"8F" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8D" , x"8D" , x"92" , x"82" , x"2F" , x"62" , x"7F" , x"7B" , x"FF" , x"A6" , x"42" , x"8D" , x"88" , x"57" , x"42" , x"51" , x"81" , x"94" , x"4B" , x"A1" , x"FE" , x"A9" , x"61" , x"7E" , x"7D" , x"75" , x"84" , x"60" , x"F7" , x"FF" , x"FE" , x"B5" , x"58" , x"88" , x"3F" , x"E7" , x"FF" , x"FD" , x"FE" , x"FF" , x"F1" , x"61" , x"81" , x"7B" , x"FF" , x"D0" , x"58" , x"79" , x"A4" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FC" , x"FF" , x"91" , x"42" , x"55" , x"51" , x"51" , x"51" , x"50" , x"51" , x"46" , x"3F" , x"83" , x"53" , x"F7" , x"F8" , x"51" , x"8B" , x"5E" , x"4F" , x"53" , x"51" , x"50" , x"50" , x"51" , x"50" , x"50" , x"50" , x"4F" , x"50" , x"50" , x"50" , x"50" , x"50" , x"4F" , x"4F" , x"4F" , x"4F" , x"4F" , x"4F" , x"4F" , x"4F" , x"4F" , x"50" , x"50" , x"50" , x"4D" , x"33" , x"72" , x"6B" , x"AA" , x"FF" , x"6A" , x"68" , x"96" , x"4B" , x"30" , x"2F" , x"31" , x"45" , x"91" , x"72" , x"67" , x"FF" , x"DA" , x"4E" , x"86" , x"54" , x"55" , x"83" , x"5E" , x"F7" , x"FF" , x"FF" , x"ED" , x"4C" , x"8C" , x"53" , x"B1" , x"FF" , x"FC" , x"FE" , x"FF" , x"F0" , x"5F" , x"81" , x"80" , x"FF" , x"CF" , x"58" , x"79" , x"A4" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FD" , x"FF" , x"E6" , x"44" , x"33" , x"31" , x"31" , x"30" , x"30" , x"32" , x"3F" , x"47" , x"83" , x"53" , x"F9" , x"F0" , x"55" , x"83" , x"37" , x"33" , x"31" , x"32" , x"31" , x"33" , x"35" , x"34" , x"33" , x"33" , x"33" , x"34" , x"3A" , x"36" , x"31" , x"33" , x"33" , x"33" , x"33" , x"33" , x"33" , x"33" , x"33" , x"33" , x"33" , x"34" , x"34" , x"33" , x"30" , x"32" , x"7E" , x"57" , x"D4" , x"FD" , x"49" , x"89" , x"70" , x"2F" , x"89" , x"C0" , x"81" , x"30" , x"64" , x"8E" , x"4A" , x"F2" , x"FC" , x"58" , x"88" , x"3E" , x"2F" , x"83" , x"5D" , x"F8" , x"FF" , x"FD" , x"FF" , x"6D" , x"7C" , x"73" , x"7B" , x"FF" , x"FC" , x"FE" , x"FF" , x"EF" , x"5F" , x"81" , x"84" , x"FF" , x"CF" , x"58" , x"79" , x"A5" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"DE" , x"B6" , x"B3" , x"AB" , x"B3" , x"B6" , x"B0" , x"D7" , x"72" , x"85" , x"57" , x"FB" , x"ED" , x"58" , x"7D" , x"5A" , x"9F" , x"9B" , x"A7" , x"AA" , x"AB" , x"94" , x"39" , x"27" , x"28" , x"34" , x"BD" , x"E7" , x"D5" , x"D2" , x"79" , x"28" , x"27" , x"26" , x"25" , x"25" , x"25" , x"25" , x"25" , x"25" , x"24" , x"24" , x"27" , x"1F" , x"33" , x"85" , x"54" , x"F7" , x"D8" , x"4B" , x"91" , x"48" , x"8C" , x"FF" , x"FF" , x"FF" , x"8F" , x"3F" , x"8E" , x"57" , x"C7" , x"FF" , x"6F" , x"83" , x"4F" , x"30" , x"82" , x"5D" , x"F7" , x"FF" , x"FB" , x"FE" , x"A6" , x"5F" , x"89" , x"52" , x"FA" , x"FF" , x"FC" , x"FD" , x"F0" , x"62" , x"81" , x"89" , x"FF" , x"CF" , x"58" , x"79" , x"A4" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7A" , x"85" , x"59" , x"FC" , x"EE" , x"5F" , x"7D" , x"A0" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"72" , x"2F" , x"2F" , x"37" , x"72" , x"A9" , x"FF" , x"FF" , x"97" , x"2F" , x"2E" , x"2E" , x"2E" , x"2E" , x"2E" , x"2E" , x"2F" , x"2E" , x"2E" , x"2E" , x"2E" , x"27" , x"42" , x"87" , x"5E" , x"FF" , x"AA" , x"69" , x"80" , x"47" , x"F5" , x"FD" , x"FB" , x"FD" , x"FB" , x"4F" , x"76" , x"74" , x"9A" , x"FF" , x"8D" , x"7A" , x"5E" , x"32" , x"82" , x"5D" , x"F6" , x"FF" , x"FD" , x"FF" , x"DE" , x"45" , x"8E" , x"4D" , x"D1" , x"FD" , x"FF" , x"FF" , x"FD" , x"64" , x"80" , x"8A" , x"FF" , x"CF" , x"58" , x"7A" , x"A5" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FD" , x"FC" , x"FC" , x"FC" , x"FC" , x"FB" , x"FD" , x"77" , x"84" , x"5A" , x"FC" , x"EE" , x"60" , x"7E" , x"A5" , x"FD" , x"F9" , x"FD" , x"FB" , x"FC" , x"D9" , x"3F" , x"3F" , x"3D" , x"3D" , x"40" , x"40" , x"C1" , x"E7" , x"39" , x"3D" , x"3F" , x"3D" , x"3D" , x"3E" , x"3C" , x"3C" , x"3C" , x"3C" , x"3B" , x"3C" , x"3B" , x"37" , x"51" , x"83" , x"71" , x"FF" , x"81" , x"7D" , x"66" , x"8F" , x"FF" , x"FC" , x"FF" , x"FC" , x"FF" , x"A4" , x"5A" , x"85" , x"7D" , x"FF" , x"AC" , x"6E" , x"6A" , x"36" , x"82" , x"5B" , x"F5" , x"FF" , x"FE" , x"FE" , x"FE" , x"5D" , x"80" , x"6B" , x"97" , x"FF" , x"DF" , x"B9" , x"92" , x"57" , x"81" , x"8C" , x"FF" , x"CF" , x"58" , x"79" , x"A5" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"78" , x"85" , x"5C" , x"FD" , x"EE" , x"5F" , x"7D" , x"A5" , x"FF" , x"FC" , x"FF" , x"FC" , x"FF" , x"95" , x"5D" , x"8A" , x"81" , x"82" , x"8A" , x"77" , x"7E" , x"9C" , x"64" , x"8A" , x"83" , x"82" , x"81" , x"80" , x"7F" , x"7F" , x"7E" , x"7D" , x"7D" , x"7B" , x"82" , x"70" , x"5A" , x"7D" , x"8B" , x"FF" , x"69" , x"86" , x"51" , x"D8" , x"FE" , x"FD" , x"FF" , x"FD" , x"FE" , x"E9" , x"50" , x"89" , x"6E" , x"FF" , x"C8" , x"64" , x"71" , x"3A" , x"81" , x"5A" , x"F3" , x"FF" , x"FE" , x"FC" , x"FF" , x"91" , x"65" , x"82" , x"67" , x"B1" , x"40" , x"32" , x"2F" , x"51" , x"7F" , x"8C" , x"FF" , x"CF" , x"58" , x"79" , x"A5" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"76" , x"85" , x"5D" , x"FE" , x"EE" , x"5E" , x"7D" , x"A6" , x"FF" , x"FC" , x"FF" , x"FC" , x"FF" , x"79" , x"80" , x"9C" , x"93" , x"94" , x"94" , x"93" , x"51" , x"44" , x"88" , x"97" , x"94" , x"95" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"94" , x"98" , x"7A" , x"62" , x"77" , x"A2" , x"FF" , x"5F" , x"89" , x"62" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"6C" , x"85" , x"63" , x"FC" , x"DD" , x"59" , x"78" , x"3B" , x"81" , x"58" , x"F1" , x"FF" , x"FE" , x"FD" , x"FF" , x"CA" , x"47" , x"8D" , x"48" , x"33" , x"45" , x"4A" , x"45" , x"5C" , x"7F" , x"89" , x"FF" , x"CF" , x"58" , x"79" , x"A5" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"75" , x"85" , x"5D" , x"FE" , x"EE" , x"5E" , x"7D" , x"A6" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"72" , x"86" , x"73" , x"6B" , x"6F" , x"6A" , x"86" , x"55" , x"43" , x"88" , x"6D" , x"6D" , x"6D" , x"6F" , x"70" , x"71" , x"73" , x"73" , x"76" , x"76" , x"73" , x"81" , x"73" , x"66" , x"70" , x"B2" , x"FD" , x"5B" , x"86" , x"7C" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"81" , x"7D" , x"5D" , x"E6" , x"EB" , x"55" , x"7C" , x"3D" , x"81" , x"55" , x"EE" , x"FF" , x"FE" , x"FE" , x"FF" , x"F5" , x"48" , x"85" , x"61" , x"47" , x"8A" , x"8B" , x"8A" , x"90" , x"80" , x"84" , x"FF" , x"CE" , x"58" , x"79" , x"A5" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"73" , x"84" , x"5D" , x"FE" , x"EC" , x"5F" , x"7D" , x"A5" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"6E" , x"83" , x"41" , x"35" , x"39" , x"31" , x"73" , x"5A" , x"4C" , x"7E" , x"36" , x"37" , x"37" , x"37" , x"36" , x"37" , x"37" , x"38" , x"39" , x"3C" , x"34" , x"60" , x"6F" , x"65" , x"6D" , x"BD" , x"EF" , x"59" , x"7E" , x"8F" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"93" , x"75" , x"60" , x"D3" , x"F6" , x"57" , x"7F" , x"3E" , x"81" , x"53" , x"ED" , x"FF" , x"FE" , x"FF" , x"FD" , x"FF" , x"77" , x"6F" , x"6E" , x"66" , x"99" , x"92" , x"92" , x"9A" , x"87" , x"83" , x"FF" , x"CD" , x"57" , x"79" , x"A4" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"73" , x"84" , x"5D" , x"FF" , x"E9" , x"5E" , x"7D" , x"A5" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"6B" , x"84" , x"45" , x"47" , x"68" , x"50" , x"78" , x"5B" , x"4B" , x"7F" , x"56" , x"5F" , x"35" , x"2B" , x"29" , x"2B" , x"36" , x"4E" , x"63" , x"7A" , x"4D" , x"71" , x"65" , x"69" , x"68" , x"C3" , x"DF" , x"5C" , x"77" , x"9E" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"9F" , x"6C" , x"68" , x"BF" , x"FD" , x"56" , x"80" , x"40" , x"80" , x"53" , x"EC" , x"FF" , x"FE" , x"FF" , x"FC" , x"FF" , x"B5" , x"64" , x"6B" , x"71" , x"72" , x"61" , x"64" , x"69" , x"60" , x"8F" , x"FF" , x"CC" , x"57" , x"79" , x"A4" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"75" , x"84" , x"5D" , x"FF" , x"E5" , x"5C" , x"7C" , x"A5" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"6D" , x"85" , x"59" , x"E9" , x"FF" , x"8D" , x"79" , x"5D" , x"4E" , x"81" , x"85" , x"FC" , x"D7" , x"C8" , x"C5" , x"CF" , x"E0" , x"F3" , x"FE" , x"FF" , x"83" , x"80" , x"5A" , x"6B" , x"64" , x"C6" , x"D7" , x"61" , x"72" , x"AB" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"AF" , x"66" , x"6D" , x"B5" , x"FF" , x"54" , x"80" , x"41" , x"80" , x"51" , x"EC" , x"FF" , x"FD" , x"FC" , x"FB" , x"FC" , x"D6" , x"66" , x"6C" , x"72" , x"50" , x"31" , x"36" , x"36" , x"37" , x"BC" , x"FF" , x"CB" , x"57" , x"79" , x"A3" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"76" , x"84" , x"5D" , x"FF" , x"E5" , x"5C" , x"7D" , x"A5" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"6E" , x"86" , x"6A" , x"FF" , x"FF" , x"93" , x"79" , x"5E" , x"4D" , x"81" , x"81" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"68" , x"8A" , x"49" , x"6F" , x"63" , x"C9" , x"D0" , x"64" , x"6E" , x"AF" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"B9" , x"61" , x"70" , x"B0" , x"FF" , x"53" , x"81" , x"41" , x"80" , x"52" , x"EC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"DF" , x"65" , x"6B" , x"75" , x"55" , x"6A" , x"71" , x"71" , x"9F" , x"FA" , x"FF" , x"CE" , x"57" , x"79" , x"A2" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"76" , x"84" , x"5C" , x"FF" , x"E4" , x"5A" , x"7D" , x"A5" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"70" , x"87" , x"68" , x"FE" , x"FF" , x"8E" , x"77" , x"5E" , x"4D" , x"81" , x"7C" , x"FE" , x"FB" , x"FD" , x"FC" , x"FC" , x"FC" , x"FB" , x"FD" , x"D1" , x"51" , x"89" , x"3A" , x"71" , x"63" , x"C7" , x"CD" , x"65" , x"6D" , x"AD" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"BD" , x"61" , x"70" , x"AF" , x"FF" , x"53" , x"80" , x"41" , x"80" , x"51" , x"EB" , x"FF" , x"F3" , x"AD" , x"A1" , x"9F" , x"6B" , x"64" , x"6D" , x"76" , x"66" , x"F7" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"CF" , x"57" , x"79" , x"A1" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"76" , x"84" , x"5C" , x"FF" , x"E4" , x"5B" , x"7E" , x"A5" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"70" , x"86" , x"68" , x"FF" , x"FF" , x"8C" , x"78" , x"5F" , x"4D" , x"81" , x"79" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"71" , x"70" , x"7E" , x"2D" , x"73" , x"62" , x"C0" , x"D1" , x"64" , x"70" , x"A8" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"B9" , x"65" , x"6F" , x"B3" , x"FF" , x"51" , x"81" , x"40" , x"80" , x"51" , x"E8" , x"FF" , x"94" , x"36" , x"32" , x"35" , x"2D" , x"62" , x"6B" , x"76" , x"6A" , x"F6" , x"FE" , x"FD" , x"FD" , x"FC" , x"FF" , x"D0" , x"58" , x"79" , x"A0" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"76" , x"84" , x"5C" , x"FF" , x"E4" , x"5B" , x"7D" , x"A6" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"71" , x"86" , x"68" , x"FF" , x"FF" , x"87" , x"78" , x"5E" , x"4A" , x"81" , x"74" , x"FF" , x"FD" , x"FF" , x"FF" , x"E4" , x"EF" , x"FF" , x"B6" , x"3D" , x"8A" , x"5F" , x"36" , x"6F" , x"67" , x"BA" , x"D9" , x"5D" , x"75" , x"9C" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"AA" , x"6B" , x"6A" , x"BA" , x"FA" , x"52" , x"81" , x"40" , x"80" , x"51" , x"E9" , x"FF" , x"64" , x"52" , x"51" , x"51" , x"48" , x"6F" , x"6A" , x"75" , x"53" , x"DA" , x"FF" , x"FD" , x"FF" , x"FD" , x"FF" , x"D0" , x"58" , x"79" , x"9F" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"76" , x"85" , x"5A" , x"FF" , x"E4" , x"5B" , x"7D" , x"A7" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"71" , x"86" , x"68" , x"FF" , x"FF" , x"82" , x"78" , x"5E" , x"4A" , x"81" , x"64" , x"FF" , x"FD" , x"FF" , x"B1" , x"40" , x"51" , x"62" , x"34" , x"5E" , x"90" , x"49" , x"7F" , x"69" , x"6C" , x"B3" , x"E6" , x"56" , x"7B" , x"8D" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"98" , x"72" , x"62" , x"C8" , x"F1" , x"53" , x"7F" , x"3E" , x"81" , x"50" , x"EB" , x"FF" , x"60" , x"8F" , x"8F" , x"8C" , x"8B" , x"94" , x"5C" , x"7B" , x"5A" , x"A0" , x"FF" , x"FC" , x"FF" , x"FD" , x"FF" , x"D1" , x"58" , x"79" , x"9E" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"75" , x"85" , x"5A" , x"FF" , x"E3" , x"5A" , x"7C" , x"A7" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"73" , x"86" , x"68" , x"FF" , x"FF" , x"80" , x"78" , x"5F" , x"49" , x"86" , x"46" , x"E7" , x"FE" , x"FF" , x"66" , x"3A" , x"35" , x"34" , x"47" , x"8E" , x"77" , x"57" , x"B7" , x"65" , x"70" , x"A5" , x"F4" , x"53" , x"83" , x"78" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"82" , x"7C" , x"5B" , x"DC" , x"E5" , x"50" , x"7D" , x"3E" , x"81" , x"50" , x"EB" , x"FF" , x"5D" , x"8D" , x"94" , x"91" , x"92" , x"90" , x"45" , x"78" , x"74" , x"5E" , x"FF" , x"FE" , x"FF" , x"FD" , x"FF" , x"D2" , x"58" , x"79" , x"9E" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"73" , x"84" , x"5A" , x"FF" , x"E3" , x"5A" , x"7C" , x"A7" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"74" , x"86" , x"68" , x"FF" , x"FF" , x"80" , x"79" , x"5F" , x"40" , x"91" , x"55" , x"9A" , x"FF" , x"FF" , x"64" , x"6E" , x"6F" , x"63" , x"85" , x"96" , x"4D" , x"8D" , x"D5" , x"5E" , x"76" , x"91" , x"FE" , x"4F" , x"89" , x"61" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"69" , x"85" , x"58" , x"F1" , x"D4" , x"58" , x"78" , x"3B" , x"81" , x"51" , x"EB" , x"FF" , x"59" , x"86" , x"60" , x"5C" , x"62" , x"54" , x"32" , x"5A" , x"89" , x"3C" , x"E2" , x"FF" , x"FD" , x"FD" , x"FF" , x"D2" , x"58" , x"79" , x"9D" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"70" , x"84" , x"5A" , x"FF" , x"E3" , x"5A" , x"7D" , x"A7" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"74" , x"86" , x"68" , x"FF" , x"FF" , x"82" , x"78" , x"5F" , x"2A" , x"7D" , x"77" , x"4B" , x"FA" , x"FF" , x"69" , x"75" , x"98" , x"91" , x"97" , x"6E" , x"33" , x"E3" , x"D9" , x"55" , x"7D" , x"7C" , x"FF" , x"52" , x"89" , x"50" , x"E4" , x"FF" , x"FD" , x"FF" , x"FE" , x"FF" , x"F1" , x"50" , x"8A" , x"57" , x"FF" , x"BE" , x"63" , x"72" , x"3A" , x"81" , x"51" , x"EB" , x"FF" , x"5A" , x"82" , x"3C" , x"32" , x"36" , x"34" , x"92" , x"4C" , x"8E" , x"52" , x"AC" , x"FF" , x"FC" , x"FD" , x"FF" , x"D2" , x"58" , x"79" , x"9D" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6F" , x"84" , x"5A" , x"FF" , x"E3" , x"5A" , x"7D" , x"A7" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"74" , x"86" , x"6A" , x"FF" , x"FF" , x"87" , x"78" , x"5D" , x"2B" , x"59" , x"8F" , x"3B" , x"C3" , x"FE" , x"8D" , x"4C" , x"90" , x"8B" , x"72" , x"3D" , x"7D" , x"FF" , x"DB" , x"50" , x"83" , x"65" , x"FF" , x"5C" , x"80" , x"5E" , x"AB" , x"FF" , x"FC" , x"FF" , x"FC" , x"FE" , x"B9" , x"54" , x"86" , x"61" , x"FF" , x"A5" , x"6D" , x"6B" , x"36" , x"81" , x"51" , x"EC" , x"FF" , x"5B" , x"84" , x"53" , x"96" , x"8E" , x"C8" , x"FF" , x"62" , x"7E" , x"6F" , x"74" , x"FF" , x"FD" , x"FD" , x"FF" , x"D2" , x"58" , x"79" , x"9C" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6F" , x"84" , x"5C" , x"FF" , x"E3" , x"5A" , x"7D" , x"A7" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"74" , x"86" , x"6B" , x"FF" , x"FF" , x"8D" , x"78" , x"5D" , x"8B" , x"45" , x"8D" , x"5A" , x"75" , x"FF" , x"CC" , x"32" , x"86" , x"6B" , x"38" , x"5F" , x"EC" , x"FF" , x"ED" , x"52" , x"87" , x"52" , x"FF" , x"73" , x"6E" , x"76" , x"5A" , x"FF" , x"FC" , x"FC" , x"FB" , x"FF" , x"63" , x"6F" , x"79" , x"7A" , x"FF" , x"89" , x"7A" , x"60" , x"31" , x"82" , x"51" , x"EC" , x"FF" , x"5E" , x"85" , x"6B" , x"FF" , x"FF" , x"FF" , x"FE" , x"9B" , x"61" , x"84" , x"49" , x"F7" , x"FF" , x"FD" , x"FF" , x"D2" , x"58" , x"79" , x"9C" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6E" , x"84" , x"5C" , x"FF" , x"E3" , x"5A" , x"7D" , x"A8" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"74" , x"86" , x"6D" , x"FF" , x"FF" , x"90" , x"77" , x"5B" , x"CB" , x"5F" , x"77" , x"7B" , x"3C" , x"EF" , x"FD" , x"4B" , x"6A" , x"83" , x"39" , x"D4" , x"FF" , x"FF" , x"FD" , x"59" , x"87" , x"46" , x"F4" , x"A4" , x"55" , x"8E" , x"3E" , x"A9" , x"FF" , x"FF" , x"FF" , x"BD" , x"38" , x"8A" , x"61" , x"A5" , x"FF" , x"67" , x"83" , x"50" , x"2E" , x"82" , x"51" , x"EC" , x"FF" , x"60" , x"86" , x"68" , x"FC" , x"FD" , x"FB" , x"FF" , x"DA" , x"47" , x"8D" , x"49" , x"CE" , x"FF" , x"FB" , x"FF" , x"D1" , x"58" , x"79" , x"9C" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6E" , x"84" , x"5D" , x"FF" , x"E2" , x"5A" , x"7D" , x"A9" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"74" , x"86" , x"6E" , x"FF" , x"FF" , x"91" , x"78" , x"5C" , x"D2" , x"AB" , x"57" , x"94" , x"41" , x"B1" , x"FF" , x"94" , x"49" , x"93" , x"4A" , x"C5" , x"FD" , x"FB" , x"FF" , x"66" , x"83" , x"53" , x"CD" , x"DD" , x"39" , x"90" , x"60" , x"32" , x"A8" , x"DA" , x"A9" , x"37" , x"57" , x"92" , x"46" , x"DF" , x"FA" , x"4C" , x"88" , x"41" , x"30" , x"82" , x"51" , x"ED" , x"FF" , x"60" , x"86" , x"64" , x"FF" , x"FF" , x"FE" , x"FE" , x"FD" , x"59" , x"82" , x"69" , x"97" , x"FF" , x"FA" , x"FF" , x"D0" , x"58" , x"79" , x"9B" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6E" , x"84" , x"5D" , x"FF" , x"E1" , x"5A" , x"7C" , x"A9" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"73" , x"86" , x"70" , x"FF" , x"FF" , x"92" , x"78" , x"5B" , x"CA" , x"F2" , x"3F" , x"8C" , x"5D" , x"70" , x"FF" , x"E3" , x"3A" , x"85" , x"6A" , x"7B" , x"FF" , x"FA" , x"FF" , x"79" , x"77" , x"68" , x"9C" , x"FF" , x"41" , x"73" , x"8C" , x"3E" , x"30" , x"36" , x"32" , x"38" , x"85" , x"7C" , x"54" , x"FF" , x"D0" , x"4A" , x"88" , x"5D" , x"5F" , x"84" , x"54" , x"ED" , x"FF" , x"60" , x"85" , x"61" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"8F" , x"67" , x"81" , x"62" , x"FF" , x"FD" , x"FF" , x"CE" , x"57" , x"79" , x"9C" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6C" , x"84" , x"5E" , x"FF" , x"E1" , x"5B" , x"7C" , x"A8" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"73" , x"87" , x"73" , x"FF" , x"FF" , x"94" , x"78" , x"5B" , x"C4" , x"FF" , x"65" , x"72" , x"7F" , x"3E" , x"EE" , x"FF" , x"6A" , x"67" , x"86" , x"42" , x"EE" , x"FE" , x"FF" , x"98" , x"64" , x"7B" , x"69" , x"FF" , x"83" , x"4D" , x"98" , x"7A" , x"42" , x"39" , x"41" , x"73" , x"9A" , x"55" , x"87" , x"FE" , x"99" , x"5F" , x"80" , x"82" , x"77" , x"84" , x"54" , x"ED" , x"FF" , x"61" , x"85" , x"61" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"CC" , x"48" , x"8E" , x"4C" , x"E4" , x"FF" , x"FF" , x"CC" , x"57" , x"79" , x"9C" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6C" , x"84" , x"60" , x"FF" , x"E1" , x"5B" , x"7C" , x"A7" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"71" , x"87" , x"74" , x"FF" , x"FF" , x"94" , x"78" , x"5A" , x"C6" , x"FE" , x"A6" , x"51" , x"95" , x"42" , x"AE" , x"FE" , x"B5" , x"45" , x"92" , x"4C" , x"A9" , x"FF" , x"FF" , x"BA" , x"4D" , x"87" , x"44" , x"F5" , x"DD" , x"31" , x"72" , x"98" , x"84" , x"74" , x"81" , x"96" , x"78" , x"37" , x"D6" , x"FF" , x"5E" , x"77" , x"6D" , x"9D" , x"77" , x"84" , x"54" , x"ED" , x"FF" , x"61" , x"85" , x"60" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F6" , x"4D" , x"87" , x"62" , x"AC" , x"FE" , x"FF" , x"C8" , x"58" , x"79" , x"9B" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6C" , x"85" , x"60" , x"FF" , x"DF" , x"59" , x"7C" , x"A8" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"71" , x"87" , x"74" , x"FF" , x"FF" , x"95" , x"78" , x"5A" , x"C9" , x"FF" , x"E5" , x"3E" , x"86" , x"63" , x"67" , x"FF" , x"F3" , x"46" , x"80" , x"6C" , x"5A" , x"FF" , x"FF" , x"DF" , x"3D" , x"8A" , x"4D" , x"B6" , x"FF" , x"67" , x"40" , x"83" , x"95" , x"92" , x"95" , x"86" , x"47" , x"65" , x"FF" , x"E0" , x"39" , x"87" , x"57" , x"C1" , x"70" , x"84" , x"56" , x"EF" , x"FF" , x"61" , x"85" , x"60" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"7D" , x"6E" , x"7D" , x"72" , x"FF" , x"FF" , x"C5" , x"58" , x"79" , x"99" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6B" , x"85" , x"60" , x"FF" , x"DF" , x"59" , x"7C" , x"A7" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"71" , x"87" , x"73" , x"FF" , x"FF" , x"97" , x"78" , x"5A" , x"CB" , x"FF" , x"FF" , x"6B" , x"6E" , x"82" , x"3A" , x"E5" , x"FF" , x"80" , x"64" , x"89" , x"39" , x"DD" , x"FF" , x"FC" , x"4F" , x"7F" , x"68" , x"69" , x"FF" , x"D7" , x"33" , x"47" , x"6E" , x"7F" , x"71" , x"4B" , x"32" , x"CD" , x"FF" , x"8F" , x"4B" , x"8C" , x"44" , x"E5" , x"68" , x"84" , x"57" , x"F1" , x"FF" , x"60" , x"85" , x"61" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"BB" , x"4F" , x"8D" , x"4D" , x"E9" , x"FF" , x"C1" , x"58" , x"79" , x"99" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6C" , x"85" , x"60" , x"FF" , x"DE" , x"59" , x"7B" , x"A7" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"71" , x"87" , x"71" , x"FF" , x"FF" , x"99" , x"78" , x"5A" , x"CC" , x"FF" , x"FF" , x"B5" , x"4D" , x"93" , x"47" , x"A8" , x"FE" , x"C2" , x"42" , x"90" , x"50" , x"9E" , x"FF" , x"FF" , x"76" , x"68" , x"84" , x"37" , x"DE" , x"FF" , x"95" , x"2F" , x"36" , x"3B" , x"37" , x"30" , x"81" , x"FF" , x"F4" , x"3E" , x"6C" , x"81" , x"50" , x"FE" , x"5D" , x"83" , x"59" , x"F2" , x"FF" , x"5E" , x"86" , x"63" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"EF" , x"47" , x"8A" , x"5B" , x"AB" , x"FE" , x"BD" , x"58" , x"79" , x"99" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6C" , x"85" , x"60" , x"FF" , x"DE" , x"59" , x"7B" , x"A8" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"71" , x"86" , x"6E" , x"FF" , x"FF" , x"99" , x"78" , x"5B" , x"CD" , x"FF" , x"FE" , x"F2" , x"48" , x"85" , x"69" , x"68" , x"FF" , x"F8" , x"4B" , x"7E" , x"71" , x"5C" , x"FE" , x"FF" , x"B1" , x"49" , x"94" , x"4E" , x"82" , x"FF" , x"FE" , x"90" , x"31" , x"2F" , x"29" , x"71" , x"F6" , x"FF" , x"A5" , x"38" , x"8D" , x"66" , x"7C" , x"FF" , x"56" , x"83" , x"56" , x"F1" , x"FF" , x"5D" , x"87" , x"65" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"73" , x"75" , x"79" , x"68" , x"FF" , x"BD" , x"58" , x"79" , x"99" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6C" , x"85" , x"5E" , x"FF" , x"DE" , x"59" , x"7B" , x"A8" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"71" , x"85" , x"6A" , x"FF" , x"FF" , x"9B" , x"78" , x"5A" , x"CD" , x"FF" , x"FA" , x"FF" , x"7C" , x"68" , x"86" , x"3B" , x"E6" , x"FF" , x"8F" , x"5F" , x"8C" , x"39" , x"D4" , x"FE" , x"E6" , x"3B" , x"84" , x"72" , x"34" , x"D4" , x"FF" , x"FF" , x"D5" , x"A9" , x"C5" , x"FF" , x"FF" , x"EF" , x"3E" , x"56" , x"93" , x"46" , x"B8" , x"FF" , x"58" , x"83" , x"55" , x"F0" , x"FF" , x"5B" , x"86" , x"67" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FE" , x"B2" , x"54" , x"8B" , x"40" , x"F4" , x"C5" , x"58" , x"79" , x"9A" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6E" , x"84" , x"5D" , x"FE" , x"DF" , x"5B" , x"7B" , x"A9" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"71" , x"86" , x"6B" , x"FD" , x"FC" , x"9C" , x"78" , x"5A" , x"CD" , x"FF" , x"FA" , x"FE" , x"C0" , x"48" , x"91" , x"4B" , x"A3" , x"FE" , x"D9" , x"43" , x"91" , x"54" , x"88" , x"FF" , x"FF" , x"63" , x"63" , x"94" , x"44" , x"59" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"7F" , x"34" , x"7F" , x"7B" , x"3B" , x"EE" , x"FF" , x"5A" , x"83" , x"53" , x"EC" , x"FE" , x"59" , x"85" , x"67" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"EA" , x"46" , x"8B" , x"54" , x"BC" , x"CE" , x"59" , x"79" , x"98" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6E" , x"85" , x"5B" , x"FF" , x"E0" , x"5A" , x"7C" , x"AA" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"71" , x"86" , x"68" , x"FF" , x"FF" , x"9E" , x"79" , x"5B" , x"CC" , x"FF" , x"FD" , x"FF" , x"F6" , x"4C" , x"83" , x"6B" , x"57" , x"FF" , x"FE" , x"5E" , x"7C" , x"73" , x"43" , x"F3" , x"FF" , x"AA" , x"3F" , x"8F" , x"70" , x"33" , x"76" , x"E4" , x"FF" , x"FF" , x"FF" , x"EC" , x"8E" , x"2C" , x"56" , x"9A" , x"59" , x"6B" , x"FF" , x"FF" , x"5D" , x"83" , x"50" , x"ED" , x"FF" , x"54" , x"85" , x"67" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6E" , x"7B" , x"73" , x"73" , x"C5" , x"58" , x"78" , x"97" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"6E" , x"82" , x"4D" , x"F4" , x"D5" , x"56" , x"7A" , x"AF" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"71" , x"84" , x"4B" , x"A2" , x"B0" , x"61" , x"78" , x"5B" , x"CD" , x"FF" , x"FD" , x"FD" , x"FF" , x"82" , x"65" , x"8A" , x"33" , x"BB" , x"FF" , x"6B" , x"5D" , x"8D" , x"39" , x"BB" , x"FF" , x"EE" , x"3C" , x"68" , x"96" , x"55" , x"31" , x"38" , x"5D" , x"65" , x"5B" , x"3C" , x"2D" , x"3F" , x"8A" , x"82" , x"37" , x"BD" , x"FF" , x"FF" , x"61" , x"83" , x"45" , x"CA" , x"DD" , x"42" , x"86" , x"67" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FE" , x"A7" , x"5C" , x"8A" , x"45" , x"79" , x"58" , x"78" , x"96" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"70" , x"81" , x"45" , x"62" , x"56" , x"5C" , x"77" , x"B7" , x"FF" , x"FC" , x"FF" , x"FE" , x"FF" , x"73" , x"84" , x"43" , x"31" , x"32" , x"32" , x"77" , x"5B" , x"D1" , x"FF" , x"FE" , x"FD" , x"FF" , x"C7" , x"43" , x"90" , x"4E" , x"37" , x"62" , x"3D" , x"46" , x"92" , x"59" , x"8A" , x"FF" , x"FF" , x"8A" , x"40" , x"8A" , x"8C" , x"4E" , x"31" , x"31" , x"32" , x"32" , x"33" , x"3F" , x"78" , x"97" , x"53" , x"53" , x"FB" , x"FE" , x"FF" , x"63" , x"82" , x"4A" , x"45" , x"47" , x"40" , x"85" , x"6A" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"DF" , x"43" , x"8E" , x"4C" , x"2B" , x"60" , x"78" , x"97" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"74" , x"84" , x"4C" , x"36" , x"32" , x"69" , x"71" , x"C2" , x"FF" , x"FD" , x"FF" , x"FE" , x"FF" , x"74" , x"82" , x"44" , x"3D" , x"3E" , x"37" , x"75" , x"5B" , x"D8" , x"FF" , x"FD" , x"FF" , x"FF" , x"F8" , x"4C" , x"80" , x"6F" , x"2F" , x"37" , x"39" , x"32" , x"74" , x"7B" , x"7A" , x"FF" , x"FD" , x"E8" , x"38" , x"5A" , x"93" , x"8A" , x"5B" , x"40" , x"3D" , x"3E" , x"4E" , x"7E" , x"9A" , x"73" , x"33" , x"C5" , x"FF" , x"FB" , x"FF" , x"69" , x"82" , x"49" , x"35" , x"36" , x"42" , x"82" , x"6E" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"5D" , x"7F" , x"6D" , x"2C" , x"5D" , x"78" , x"9B" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"7D" , x"7D" , x"7C" , x"6D" , x"6B" , x"84" , x"62" , x"D3" , x"FF" , x"FD" , x"FF" , x"FD" , x"FF" , x"79" , x"85" , x"7E" , x"78" , x"78" , x"78" , x"8B" , x"5A" , x"E4" , x"FF" , x"FD" , x"FF" , x"FD" , x"FF" , x"84" , x"60" , x"8E" , x"6C" , x"72" , x"6E" , x"6A" , x"7F" , x"7F" , x"7F" , x"FF" , x"FA" , x"FF" , x"9F" , x"36" , x"6B" , x"93" , x"8E" , x"80" , x"77" , x"7B" , x"8A" , x"95" , x"80" , x"40" , x"74" , x"FF" , x"FE" , x"FD" , x"FF" , x"76" , x"80" , x"7A" , x"6D" , x"6D" , x"76" , x"85" , x"75" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"96" , x"61" , x"8E" , x"69" , x"82" , x"71" , x"A4" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"90" , x"6E" , x"9D" , x"93" , x"93" , x"92" , x"58" , x"EC" , x"FF" , x"FE" , x"FF" , x"FC" , x"FF" , x"85" , x"7F" , x"9C" , x"93" , x"96" , x"97" , x"92" , x"5C" , x"F7" , x"FF" , x"FE" , x"FF" , x"FD" , x"FF" , x"CC" , x"43" , x"8C" , x"95" , x"92" , x"93" , x"95" , x"9B" , x"7F" , x"85" , x"FF" , x"FB" , x"FD" , x"FA" , x"5E" , x"3C" , x"6B" , x"91" , x"95" , x"95" , x"94" , x"94" , x"7D" , x"44" , x"47" , x"EA" , x"FE" , x"FD" , x"FC" , x"FF" , x"89" , x"74" , x"9D" , x"93" , x"93" , x"9C" , x"7E" , x"81" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"D3" , x"46" , x"90" , x"94" , x"9A" , x"61" , x"B6" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"B9" , x"4D" , x"85" , x"80" , x"87" , x"76" , x"64" , x"FF" , x"FE" , x"FF" , x"FF" , x"FC" , x"FF" , x"A6" , x"54" , x"81" , x"79" , x"79" , x"80" , x"6C" , x"6B" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FE" , x"FC" , x"55" , x"75" , x"8A" , x"80" , x"83" , x"82" , x"88" , x"78" , x"95" , x"FF" , x"FC" , x"FD" , x"FF" , x"E4" , x"47" , x"38" , x"55" , x"70" , x"7A" , x"76" , x"61" , x"3E" , x"39" , x"C9" , x"FF" , x"FE" , x"FF" , x"FC" , x"FF" , x"AD" , x"50" , x"86" , x"80" , x"81" , x"88" , x"57" , x"A4" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FB" , x"56" , x"77" , x"87" , x"7D" , x"44" , x"E0" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"ED" , x"3F" , x"40" , x"43" , x"41" , x"3E" , x"AB" , x"FF" , x"FD" , x"FF" , x"FF" , x"FD" , x"FF" , x"E3" , x"39" , x"3B" , x"3A" , x"39" , x"3A" , x"3B" , x"B5" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"9B" , x"40" , x"48" , x"43" , x"43" , x"41" , x"42" , x"42" , x"B7" , x"FF" , x"FC" , x"FF" , x"FD" , x"FF" , x"D5" , x"50" , x"33" , x"35" , x"3A" , x"38" , x"33" , x"47" , x"C1" , x"FF" , x"FC" , x"FF" , x"FF" , x"FD" , x"FF" , x"E4" , x"37" , x"41" , x"44" , x"43" , x"3F" , x"3D" , x"E5" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"9B" , x"3E" , x"47" , x"3E" , x"69" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"AB" , x"34" , x"34" , x"38" , x"7B" , x"FA" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"B3" , x"55" , x"46" , x"46" , x"51" , x"98" , x"FE" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FD" , x"FE" , x"EB" , x"43" , x"35" , x"32" , x"35" , x"34" , x"37" , x"50" , x"ED" , x"FF" , x"FE" , x"FF" , x"FF" , x"FD" , x"FF" , x"EE" , x"8B" , x"4B" , x"41" , x"4B" , x"88" , x"E5" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"8D" , x"34" , x"33" , x"34" , x"35" , x"AA" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FE" , x"EE" , x"51" , x"38" , x"40" , x"D8" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"CE" , x"B7" , x"D2" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F8" , x"EA" , x"EB" , x"F6" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"CE" , x"82" , x"8D" , x"9B" , x"A1" , x"A9" , x"E3" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"FF" , x"F3" , x"E4" , x"F2" , x"FF" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FF" , x"B2" , x"8E" , x"97" , x"C7" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"E4" , x"97" , x"D3" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"FF" , x"FF" , x"FF" , x"FD" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FC" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FC" , x"FC" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FC" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ) 
);

CONSTANT Plantilla_TronG : ImageMatrix(0 TO 99, 0 TO 99) := (
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"65" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"65" , x"65" , x"64" , x"64" , x"65" , x"65" , x"66" , x"65" , x"65" , x"66" , x"65" , x"66" , x"66" , x"66" , x"65" , x"64" , x"64" , x"63" , x"64" , x"65" , x"64" , x"64" , x"66" , x"66" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"63" , x"61" , x"63" , x"63" , x"63" , x"65" , x"63" , x"64" , x"66" , x"66" , x"65" , x"62" , x"65" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"63" , x"64" , x"63" , x"63" , x"63" , x"63" , x"63" , x"62" , x"62" , x"62" , x"63" , x"63" , x"63" , x"65" , x"63" , x"61" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"61" , x"64" , x"62" , x"5E" , x"62" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"65" , x"66" , x"62" , x"64" , x"64" , x"61" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"64" , x"5A" , x"62" , x"60" , x"61" , x"60" , x"62" , x"66" , x"65" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"5C" , x"77" , x"87" , x"85" , x"86" , x"87" , x"87" , x"87" , x"86" , x"63" , x"66" , x"63" , x"60" , x"7E" , x"86" , x"86" , x"86" , x"86" , x"86" , x"86" , x"87" , x"87" , x"87" , x"87" , x"87" , x"87" , x"86" , x"87" , x"87" , x"87" , x"87" , x"87" , x"86" , x"87" , x"87" , x"86" , x"86" , x"86" , x"86" , x"82" , x"73" , x"60" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"65" , x"66" , x"61" , x"60" , x"70" , x"7F" , x"87" , x"83" , x"78" , x"64" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"65" , x"67" , x"87" , x"86" , x"7B" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"65" , x"66" , x"5A" , x"77" , x"86" , x"86" , x"85" , x"86" , x"62" , x"65" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"67" , x"66" , x"5D" , x"AF" , x"D2" , x"CD" , x"CF" , x"CF" , x"CE" , x"D0" , x"C8" , x"73" , x"63" , x"5E" , x"80" , x"B4" , x"CD" , x"CE" , x"CE" , x"CE" , x"CE" , x"CE" , x"CE" , x"CE" , x"CF" , x"CE" , x"CE" , x"CF" , x"CE" , x"CE" , x"CF" , x"CF" , x"CF" , x"CE" , x"CE" , x"CF" , x"CF" , x"CE" , x"CE" , x"CD" , x"CF" , x"C7" , x"A2" , x"80" , x"5E" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"63" , x"61" , x"82" , x"9E" , x"C3" , x"CE" , x"CA" , x"AC" , x"89" , x"68" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"66" , x"61" , x"8C" , x"CA" , x"D2" , x"BC" , x"65" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"60" , x"AF" , x"D0" , x"CD" , x"CF" , x"C7" , x"7C" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"67" , x"66" , x"6B" , x"E9" , x"FE" , x"FB" , x"FC" , x"FB" , x"FC" , x"FB" , x"FE" , x"9B" , x"58" , x"68" , x"BA" , x"F9" , x"F9" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FC" , x"FB" , x"FB" , x"FC" , x"F1" , x"B5" , x"75" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5E" , x"84" , x"BB" , x"F0" , x"FC" , x"FC" , x"FC" , x"F6" , x"D0" , x"90" , x"62" , x"62" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"C2" , x"FD" , x"FC" , x"ED" , x"77" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"73" , x"EC" , x"FE" , x"FB" , x"FB" , x"FD" , x"AC" , x"5C" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"64" , x"7B" , x"F3" , x"E5" , x"E4" , x"E3" , x"E4" , x"E5" , x"E1" , x"F4" , x"B3" , x"50" , x"8A" , x"F2" , x"F4" , x"E1" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E5" , x"E4" , x"E3" , x"E9" , x"F9" , x"F5" , x"A8" , x"61" , x"66" , x"66" , x"66" , x"66" , x"66" , x"61" , x"76" , x"C0" , x"FB" , x"FA" , x"EC" , x"E4" , x"E8" , x"F6" , x"FE" , x"D8" , x"89" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"68" , x"E0" , x"EE" , x"E1" , x"F5" , x"9E" , x"60" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"63" , x"88" , x"F7" , x"E3" , x"E4" , x"E1" , x"F1" , x"CC" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"62" , x"82" , x"EA" , x"98" , x"91" , x"92" , x"92" , x"94" , x"8B" , x"CE" , x"BF" , x"5E" , x"BC" , x"FB" , x"B0" , x"8E" , x"91" , x"91" , x"90" , x"91" , x"90" , x"92" , x"92" , x"91" , x"91" , x"92" , x"91" , x"91" , x"91" , x"91" , x"91" , x"91" , x"90" , x"91" , x"90" , x"91" , x"91" , x"90" , x"91" , x"91" , x"96" , x"BE" , x"F9" , x"E1" , x"7B" , x"61" , x"66" , x"66" , x"67" , x"65" , x"65" , x"AC" , x"F8" , x"F4" , x"C1" , x"99" , x"91" , x"94" , x"B1" , x"E5" , x"FE" , x"C8" , x"72" , x"62" , x"66" , x"67" , x"66" , x"6F" , x"E5" , x"AB" , x"8B" , x"E1" , x"CE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"62" , x"94" , x"E7" , x"91" , x"95" , x"8D" , x"B9" , x"D5" , x"62" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"62" , x"83" , x"EA" , x"85" , x"67" , x"69" , x"68" , x"6B" , x"6C" , x"CB" , x"C3" , x"79" , x"E6" , x"D0" , x"78" , x"6B" , x"69" , x"6A" , x"6A" , x"6A" , x"6A" , x"6B" , x"6B" , x"6B" , x"6B" , x"6B" , x"6A" , x"6A" , x"6A" , x"6B" , x"6B" , x"6B" , x"6A" , x"69" , x"69" , x"69" , x"69" , x"69" , x"6A" , x"6A" , x"6F" , x"7E" , x"BC" , x"FD" , x"AF" , x"60" , x"66" , x"66" , x"66" , x"5D" , x"89" , x"E8" , x"F7" , x"AB" , x"81" , x"73" , x"6A" , x"6F" , x"7C" , x"97" , x"E3" , x"FA" , x"A9" , x"61" , x"66" , x"68" , x"66" , x"73" , x"EA" , x"99" , x"68" , x"BC" , x"EE" , x"71" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"61" , x"96" , x"E4" , x"79" , x"6C" , x"6C" , x"B0" , x"DA" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"62" , x"82" , x"EF" , x"79" , x"5E" , x"60" , x"61" , x"64" , x"60" , x"CC" , x"C2" , x"92" , x"F2" , x"9E" , x"5F" , x"5D" , x"60" , x"5E" , x"5E" , x"5D" , x"5C" , x"5B" , x"59" , x"59" , x"5A" , x"5C" , x"5C" , x"5C" , x"5B" , x"5A" , x"59" , x"5A" , x"5C" , x"5D" , x"5F" , x"5E" , x"5D" , x"5D" , x"5C" , x"5C" , x"5C" , x"62" , x"80" , x"E2" , x"DF" , x"69" , x"66" , x"67" , x"64" , x"60" , x"BE" , x"FD" , x"B5" , x"75" , x"62" , x"5A" , x"5A" , x"5A" , x"5F" , x"6D" , x"9A" , x"F2" , x"E0" , x"75" , x"62" , x"66" , x"66" , x"72" , x"EE" , x"91" , x"5A" , x"92" , x"F8" , x"93" , x"60" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"96" , x"E9" , x"6C" , x"64" , x"5E" , x"B0" , x"DE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"61" , x"82" , x"F2" , x"77" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"C9" , x"BF" , x"A9" , x"ED" , x"75" , x"65" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"65" , x"62" , x"B0" , x"F5" , x"82" , x"5F" , x"66" , x"5D" , x"87" , x"F0" , x"D8" , x"7D" , x"60" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"6E" , x"B7" , x"FC" , x"AB" , x"62" , x"66" , x"66" , x"71" , x"EE" , x"8D" , x"66" , x"72" , x"EC" , x"C2" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"96" , x"EA" , x"6A" , x"66" , x"5F" , x"AB" , x"DF" , x"62" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"61" , x"82" , x"F1" , x"76" , x"66" , x"67" , x"66" , x"66" , x"5F" , x"CA" , x"BE" , x"BF" , x"DA" , x"65" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"61" , x"80" , x"F0" , x"A6" , x"5B" , x"66" , x"5C" , x"B9" , x"FB" , x"A0" , x"61" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5E" , x"84" , x"E6" , x"DC" , x"6D" , x"64" , x"66" , x"71" , x"EF" , x"8B" , x"67" , x"62" , x"CA" , x"E6" , x"6B" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"96" , x"EA" , x"69" , x"66" , x"5F" , x"AB" , x"DF" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"61" , x"82" , x"F1" , x"76" , x"66" , x"67" , x"66" , x"66" , x"5F" , x"C9" , x"BE" , x"CD" , x"C0" , x"5E" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"67" , x"67" , x"66" , x"67" , x"67" , x"66" , x"67" , x"67" , x"67" , x"67" , x"66" , x"66" , x"DC" , x"C5" , x"5B" , x"62" , x"68" , x"E4" , x"D7" , x"70" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"65" , x"61" , x"B5" , x"F7" , x"8B" , x"5E" , x"66" , x"71" , x"EF" , x"8A" , x"66" , x"60" , x"9C" , x"F5" , x"89" , x"5E" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"96" , x"EA" , x"68" , x"66" , x"5D" , x"AB" , x"DF" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"61" , x"82" , x"F1" , x"77" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"C8" , x"C1" , x"D6" , x"A7" , x"5D" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"61" , x"C3" , x"D9" , x"60" , x"59" , x"92" , x"F8" , x"A7" , x"5E" , x"66" , x"66" , x"60" , x"5B" , x"5D" , x"5C" , x"60" , x"66" , x"66" , x"5E" , x"83" , x"F1" , x"BE" , x"5C" , x"66" , x"72" , x"EF" , x"8B" , x"64" , x"64" , x"77" , x"EE" , x"BA" , x"5D" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"61" , x"96" , x"EA" , x"68" , x"66" , x"5E" , x"AA" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"61" , x"83" , x"ED" , x"7F" , x"5A" , x"5B" , x"5D" , x"5F" , x"61" , x"CB" , x"C3" , x"DC" , x"95" , x"5D" , x"66" , x"66" , x"61" , x"5D" , x"5D" , x"5B" , x"5B" , x"5A" , x"5A" , x"5A" , x"59" , x"5C" , x"5F" , x"5D" , x"5B" , x"5A" , x"58" , x"59" , x"59" , x"59" , x"5B" , x"5C" , x"59" , x"57" , x"58" , x"58" , x"59" , x"5C" , x"60" , x"64" , x"B1" , x"E4" , x"64" , x"58" , x"C1" , x"ED" , x"78" , x"61" , x"66" , x"5D" , x"60" , x"7A" , x"7E" , x"7D" , x"65" , x"5F" , x"66" , x"65" , x"61" , x"D0" , x"E4" , x"68" , x"66" , x"71" , x"EF" , x"8C" , x"61" , x"66" , x"64" , x"D1" , x"E0" , x"68" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"61" , x"96" , x"EA" , x"68" , x"66" , x"5D" , x"AA" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"62" , x"84" , x"E9" , x"89" , x"7A" , x"7B" , x"7C" , x"7B" , x"79" , x"C7" , x"C5" , x"DF" , x"8B" , x"5E" , x"66" , x"63" , x"5E" , x"7C" , x"7C" , x"7C" , x"7C" , x"7B" , x"7C" , x"7C" , x"7C" , x"7C" , x"7C" , x"7B" , x"7C" , x"7C" , x"7C" , x"7C" , x"7C" , x"7C" , x"7B" , x"7B" , x"7B" , x"7B" , x"7B" , x"7C" , x"7B" , x"7B" , x"7C" , x"7B" , x"A2" , x"E7" , x"61" , x"5E" , x"E1" , x"CD" , x"62" , x"66" , x"60" , x"5F" , x"8A" , x"AF" , x"C2" , x"B2" , x"8E" , x"64" , x"62" , x"66" , x"5D" , x"A3" , x"F4" , x"81" , x"5E" , x"74" , x"EF" , x"8B" , x"61" , x"66" , x"5D" , x"A4" , x"F4" , x"83" , x"60" , x"66" , x"66" , x"66" , x"66" , x"66" , x"61" , x"96" , x"EA" , x"67" , x"66" , x"5E" , x"AB" , x"DF" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"62" , x"81" , x"ED" , x"B3" , x"B0" , x"B1" , x"B1" , x"B3" , x"AC" , x"D9" , x"C3" , x"E0" , x"86" , x"5E" , x"66" , x"5B" , x"81" , x"AF" , x"B2" , x"B2" , x"B2" , x"B1" , x"B2" , x"B2" , x"B2" , x"B2" , x"B2" , x"B1" , x"B2" , x"B2" , x"B2" , x"B2" , x"B2" , x"B2" , x"B2" , x"B2" , x"B2" , x"B2" , x"B2" , x"B2" , x"B2" , x"B2" , x"B3" , x"AF" , x"BF" , x"E5" , x"64" , x"75" , x"F2" , x"A2" , x"5E" , x"66" , x"57" , x"85" , x"CD" , x"F8" , x"FB" , x"FA" , x"D4" , x"8B" , x"5D" , x"66" , x"62" , x"78" , x"F1" , x"A6" , x"58" , x"75" , x"F0" , x"8B" , x"62" , x"66" , x"62" , x"7B" , x"F2" , x"B0" , x"5C" , x"66" , x"66" , x"66" , x"66" , x"66" , x"61" , x"96" , x"EA" , x"67" , x"66" , x"5E" , x"AB" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"65" , x"74" , x"F2" , x"FA" , x"F8" , x"F9" , x"F9" , x"F9" , x"F8" , x"FB" , x"B8" , x"E2" , x"85" , x"5F" , x"66" , x"5B" , x"BA" , x"FA" , x"F7" , x"F9" , x"F9" , x"F9" , x"F8" , x"F7" , x"F7" , x"F6" , x"F6" , x"F6" , x"F6" , x"F6" , x"F8" , x"F9" , x"F7" , x"F6" , x"F7" , x"F8" , x"F7" , x"F7" , x"F7" , x"F7" , x"F7" , x"F7" , x"F8" , x"F8" , x"FA" , x"E6" , x"6F" , x"98" , x"F4" , x"7B" , x"65" , x"61" , x"63" , x"BE" , x"FC" , x"F5" , x"EA" , x"F3" , x"FE" , x"C9" , x"6B" , x"62" , x"66" , x"64" , x"DD" , x"CA" , x"5A" , x"73" , x"F1" , x"8C" , x"63" , x"67" , x"66" , x"65" , x"DA" , x"D9" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"61" , x"96" , x"EA" , x"67" , x"66" , x"5D" , x"AA" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"67" , x"66" , x"64" , x"D6" , x"F9" , x"F3" , x"F4" , x"F4" , x"F3" , x"F5" , x"ED" , x"A1" , x"E6" , x"84" , x"61" , x"66" , x"6A" , x"E6" , x"FA" , x"F5" , x"F5" , x"F5" , x"F5" , x"F5" , x"F6" , x"F4" , x"F3" , x"F3" , x"F3" , x"F2" , x"F3" , x"F4" , x"F4" , x"F4" , x"F3" , x"F4" , x"F4" , x"F4" , x"F4" , x"F4" , x"F4" , x"F4" , x"F4" , x"F5" , x"F5" , x"F9" , x"E4" , x"76" , x"B8" , x"E5" , x"69" , x"66" , x"5A" , x"8F" , x"F2" , x"EC" , x"AE" , x"94" , x"A9" , x"E5" , x"F9" , x"9D" , x"5D" , x"66" , x"5E" , x"BD" , x"E4" , x"61" , x"72" , x"F1" , x"8C" , x"63" , x"67" , x"66" , x"5F" , x"B0" , x"F2" , x"7B" , x"60" , x"66" , x"66" , x"66" , x"66" , x"60" , x"96" , x"EA" , x"67" , x"66" , x"5E" , x"AA" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"5E" , x"94" , x"AA" , x"A6" , x"A6" , x"A6" , x"A7" , x"A9" , x"9F" , x"90" , x"E9" , x"84" , x"63" , x"63" , x"7D" , x"F2" , x"B5" , x"A3" , x"A6" , x"A7" , x"A7" , x"A7" , x"A7" , x"A7" , x"A7" , x"A7" , x"A7" , x"A8" , x"A8" , x"A8" , x"A8" , x"A7" , x"A7" , x"A7" , x"A7" , x"A7" , x"A7" , x"A7" , x"A7" , x"A7" , x"A7" , x"A6" , x"A6" , x"A9" , x"A0" , x"7B" , x"D1" , x"CB" , x"61" , x"66" , x"60" , x"C6" , x"FB" , x"A3" , x"76" , x"6E" , x"78" , x"99" , x"F5" , x"D5" , x"67" , x"66" , x"5E" , x"98" , x"F1" , x"6E" , x"6E" , x"EF" , x"8B" , x"63" , x"66" , x"66" , x"62" , x"82" , x"F5" , x"A7" , x"5C" , x"66" , x"65" , x"66" , x"66" , x"60" , x"95" , x"EA" , x"68" , x"66" , x"5E" , x"AA" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"62" , x"66" , x"78" , x"74" , x"76" , x"75" , x"76" , x"77" , x"6C" , x"83" , x"EC" , x"84" , x"64" , x"60" , x"8F" , x"EA" , x"81" , x"74" , x"77" , x"77" , x"77" , x"76" , x"75" , x"76" , x"76" , x"76" , x"78" , x"75" , x"73" , x"73" , x"73" , x"78" , x"77" , x"76" , x"76" , x"76" , x"76" , x"76" , x"76" , x"76" , x"76" , x"76" , x"76" , x"78" , x"71" , x"77" , x"E4" , x"A9" , x"5E" , x"65" , x"75" , x"F1" , x"CD" , x"70" , x"5F" , x"5F" , x"5D" , x"6B" , x"BF" , x"F7" , x"81" , x"63" , x"65" , x"7F" , x"F4" , x"83" , x"6B" , x"EC" , x"8C" , x"63" , x"66" , x"67" , x"66" , x"68" , x"E0" , x"D2" , x"62" , x"66" , x"66" , x"66" , x"66" , x"60" , x"96" , x"EA" , x"69" , x"66" , x"5E" , x"AA" , x"DF" , x"65" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"62" , x"61" , x"60" , x"60" , x"60" , x"60" , x"62" , x"61" , x"79" , x"F1" , x"84" , x"64" , x"5F" , x"96" , x"E6" , x"6C" , x"5D" , x"5E" , x"5F" , x"60" , x"60" , x"5C" , x"57" , x"5E" , x"5D" , x"5D" , x"62" , x"64" , x"64" , x"63" , x"5D" , x"5D" , x"5D" , x"5D" , x"5E" , x"5E" , x"5E" , x"5E" , x"5E" , x"5E" , x"5E" , x"5E" , x"5F" , x"55" , x"76" , x"EE" , x"8E" , x"63" , x"5E" , x"99" , x"F7" , x"9A" , x"5E" , x"66" , x"66" , x"66" , x"5B" , x"8B" , x"F4" , x"AC" , x"60" , x"66" , x"6E" , x"EE" , x"9B" , x"71" , x"EB" , x"8B" , x"63" , x"66" , x"66" , x"66" , x"60" , x"BA" , x"EF" , x"74" , x"64" , x"66" , x"66" , x"66" , x"61" , x"96" , x"EB" , x"6A" , x"66" , x"5E" , x"AA" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"77" , x"F1" , x"84" , x"65" , x"5F" , x"98" , x"E5" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"62" , x"6E" , x"69" , x"69" , x"6B" , x"69" , x"66" , x"66" , x"65" , x"6B" , x"6A" , x"69" , x"6A" , x"6A" , x"6A" , x"69" , x"6A" , x"6A" , x"6B" , x"6A" , x"6B" , x"63" , x"8C" , x"F0" , x"7C" , x"66" , x"5E" , x"C4" , x"E3" , x"6F" , x"64" , x"66" , x"66" , x"66" , x"64" , x"64" , x"D8" , x"D5" , x"64" , x"66" , x"64" , x"E0" , x"B0" , x"78" , x"EA" , x"8A" , x"62" , x"66" , x"66" , x"66" , x"5F" , x"8A" , x"F7" , x"9A" , x"5F" , x"66" , x"66" , x"66" , x"65" , x"98" , x"EB" , x"6A" , x"66" , x"5E" , x"AA" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"76" , x"F1" , x"84" , x"65" , x"5F" , x"99" , x"E7" , x"68" , x"66" , x"66" , x"66" , x"66" , x"66" , x"63" , x"7A" , x"92" , x"8F" , x"8F" , x"95" , x"90" , x"6A" , x"65" , x"81" , x"90" , x"8D" , x"8E" , x"8D" , x"8C" , x"8B" , x"8B" , x"8C" , x"8B" , x"8A" , x"8A" , x"8D" , x"85" , x"A2" , x"EB" , x"71" , x"66" , x"65" , x"E2" , x"C4" , x"61" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5B" , x"B1" , x"ED" , x"70" , x"66" , x"60" , x"CF" , x"C2" , x"80" , x"E9" , x"8A" , x"62" , x"66" , x"66" , x"67" , x"66" , x"6D" , x"E6" , x"C9" , x"62" , x"66" , x"63" , x"5F" , x"55" , x"9B" , x"E8" , x"69" , x"66" , x"5E" , x"AA" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"76" , x"F2" , x"84" , x"65" , x"5F" , x"99" , x"E6" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"B9" , x"EB" , x"E6" , x"E5" , x"EA" , x"DA" , x"75" , x"66" , x"C5" , x"E9" , x"E4" , x"E4" , x"E4" , x"E4" , x"E3" , x"E3" , x"E2" , x"E1" , x"E1" , x"DF" , x"E4" , x"CE" , x"B1" , x"E4" , x"69" , x"66" , x"74" , x"F2" , x"9B" , x"5E" , x"66" , x"66" , x"66" , x"65" , x"66" , x"60" , x"89" , x"F6" , x"81" , x"66" , x"5D" , x"BD" , x"CF" , x"86" , x"E9" , x"8B" , x"61" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"C3" , x"EB" , x"74" , x"64" , x"6D" , x"71" , x"6D" , x"A3" , x"E6" , x"69" , x"66" , x"5E" , x"AA" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"76" , x"F2" , x"85" , x"66" , x"5F" , x"99" , x"E6" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"69" , x"E6" , x"FD" , x"FB" , x"FC" , x"FB" , x"FD" , x"90" , x"78" , x"F1" , x"FE" , x"FB" , x"FC" , x"FD" , x"FD" , x"FC" , x"FD" , x"FD" , x"FC" , x"FD" , x"FC" , x"FF" , x"DB" , x"BA" , x"DA" , x"63" , x"66" , x"85" , x"F5" , x"80" , x"65" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"73" , x"F3" , x"93" , x"65" , x"5E" , x"AB" , x"DA" , x"8A" , x"E8" , x"8A" , x"60" , x"66" , x"66" , x"66" , x"66" , x"5E" , x"94" , x"F6" , x"96" , x"77" , x"9B" , x"9F" , x"98" , x"B6" , x"E6" , x"6C" , x"66" , x"5D" , x"AB" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F2" , x"85" , x"66" , x"5F" , x"9A" , x"E6" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"77" , x"EF" , x"D0" , x"CB" , x"CF" , x"CA" , x"ED" , x"AB" , x"96" , x"EF" , x"CE" , x"CD" , x"CF" , x"CE" , x"CF" , x"D0" , x"D1" , x"D1" , x"D2" , x"D3" , x"D0" , x"E4" , x"D2" , x"BF" , x"D1" , x"62" , x"65" , x"95" , x"EF" , x"70" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"E7" , x"A6" , x"5E" , x"5E" , x"A0" , x"E0" , x"8C" , x"E7" , x"8B" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"64" , x"72" , x"EC" , x"BC" , x"9D" , x"EE" , x"EF" , x"ED" , x"F3" , x"E8" , x"6F" , x"66" , x"5D" , x"AA" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"85" , x"66" , x"5E" , x"9A" , x"E5" , x"67" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7C" , x"EC" , x"91" , x"83" , x"87" , x"81" , x"D5" , x"B3" , x"A0" , x"E0" , x"87" , x"84" , x"84" , x"83" , x"83" , x"83" , x"85" , x"85" , x"86" , x"8C" , x"85" , x"BD" , x"CC" , x"C2" , x"CA" , x"60" , x"60" , x"A4" , x"E5" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"D8" , x"B6" , x"5E" , x"62" , x"98" , x"E3" , x"8E" , x"E7" , x"8B" , x"5F" , x"66" , x"66" , x"66" , x"67" , x"66" , x"60" , x"D0" , x"C9" , x"C2" , x"FF" , x"F8" , x"FA" , x"FD" , x"ED" , x"6F" , x"66" , x"5D" , x"AB" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"85" , x"66" , x"5D" , x"9C" , x"E5" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7B" , x"EF" , x"8A" , x"5D" , x"62" , x"6D" , x"DB" , x"B2" , x"9F" , x"E5" , x"79" , x"60" , x"5D" , x"5A" , x"5A" , x"5A" , x"5C" , x"5E" , x"62" , x"68" , x"76" , x"D6" , x"BF" , x"C5" , x"C4" , x"5E" , x"5C" , x"B0" , x"DA" , x"61" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5A" , x"CC" , x"C3" , x"5D" , x"65" , x"92" , x"E5" , x"90" , x"E7" , x"8B" , x"5E" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"C0" , x"C9" , x"D1" , x"D4" , x"BB" , x"BE" , x"BF" , x"BB" , x"6B" , x"66" , x"5D" , x"AB" , x"DF" , x"65" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"76" , x"F1" , x"85" , x"66" , x"5D" , x"9F" , x"E4" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7C" , x"F2" , x"7D" , x"5F" , x"66" , x"61" , x"DC" , x"B3" , x"9F" , x"E9" , x"6F" , x"65" , x"5F" , x"5A" , x"5A" , x"5B" , x"5E" , x"62" , x"66" , x"66" , x"71" , x"EA" , x"AE" , x"C8" , x"BE" , x"5C" , x"5D" , x"BA" , x"D2" , x"5D" , x"66" , x"66" , x"66" , x"66" , x"66" , x"65" , x"66" , x"5A" , x"C2" , x"CD" , x"5F" , x"66" , x"8D" , x"E6" , x"90" , x"E6" , x"8B" , x"5E" , x"66" , x"65" , x"66" , x"66" , x"66" , x"5E" , x"BA" , x"CC" , x"D3" , x"A7" , x"81" , x"87" , x"86" , x"7D" , x"64" , x"66" , x"5C" , x"AB" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"85" , x"66" , x"5E" , x"A2" , x"E4" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7C" , x"F2" , x"7E" , x"66" , x"66" , x"61" , x"DB" , x"B3" , x"9E" , x"E9" , x"6D" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"65" , x"80" , x"F3" , x"9A" , x"CC" , x"BB" , x"5C" , x"5D" , x"BF" , x"CB" , x"5B" , x"66" , x"65" , x"66" , x"66" , x"66" , x"66" , x"66" , x"59" , x"BC" , x"D1" , x"60" , x"66" , x"8A" , x"E8" , x"91" , x"E6" , x"8B" , x"5E" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"BA" , x"CC" , x"D7" , x"A5" , x"63" , x"67" , x"68" , x"63" , x"65" , x"66" , x"5C" , x"AB" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"76" , x"F1" , x"84" , x"66" , x"5E" , x"A2" , x"E4" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7C" , x"F2" , x"7E" , x"66" , x"66" , x"5F" , x"DC" , x"B3" , x"9E" , x"E9" , x"6E" , x"66" , x"67" , x"66" , x"66" , x"65" , x"66" , x"66" , x"66" , x"60" , x"A4" , x"ED" , x"8A" , x"CF" , x"BB" , x"5B" , x"5C" , x"BF" , x"CB" , x"5B" , x"66" , x"65" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5A" , x"BB" , x"D0" , x"60" , x"66" , x"8A" , x"E8" , x"90" , x"E6" , x"8B" , x"5E" , x"66" , x"64" , x"5F" , x"5F" , x"5D" , x"5B" , x"C0" , x"CB" , x"DA" , x"9F" , x"63" , x"66" , x"66" , x"66" , x"67" , x"66" , x"5D" , x"AB" , x"DF" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"76" , x"F1" , x"84" , x"66" , x"5E" , x"A1" , x"E4" , x"67" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7C" , x"F2" , x"7E" , x"66" , x"66" , x"60" , x"DB" , x"B3" , x"9E" , x"E9" , x"6C" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"64" , x"D4" , x"DA" , x"78" , x"CF" , x"BE" , x"5B" , x"5C" , x"BC" , x"CF" , x"5C" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5B" , x"BF" , x"CE" , x"5F" , x"66" , x"8D" , x"E6" , x"91" , x"E6" , x"8A" , x"5D" , x"66" , x"65" , x"78" , x"75" , x"75" , x"75" , x"BD" , x"C7" , x"DB" , x"9D" , x"62" , x"67" , x"66" , x"66" , x"66" , x"66" , x"5D" , x"AB" , x"DE" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"76" , x"F1" , x"84" , x"66" , x"5E" , x"A1" , x"E4" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F2" , x"7E" , x"66" , x"66" , x"5F" , x"DB" , x"B3" , x"9D" , x"E9" , x"6D" , x"66" , x"67" , x"66" , x"66" , x"5F" , x"62" , x"66" , x"60" , x"84" , x"F0" , x"B6" , x"5F" , x"CB" , x"C4" , x"5C" , x"5C" , x"B4" , x"D7" , x"5E" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5B" , x"C8" , x"C7" , x"5E" , x"64" , x"92" , x"E5" , x"90" , x"E7" , x"8A" , x"5D" , x"66" , x"74" , x"A9" , x"A3" , x"A3" , x"9E" , x"CF" , x"C4" , x"D8" , x"9F" , x"5E" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5C" , x"AB" , x"DE" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"84" , x"66" , x"5E" , x"A2" , x"E4" , x"67" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F2" , x"7E" , x"66" , x"66" , x"5E" , x"DB" , x"B4" , x"9C" , x"E8" , x"72" , x"66" , x"67" , x"66" , x"5B" , x"5E" , x"5F" , x"5F" , x"6C" , x"BC" , x"F9" , x"8A" , x"57" , x"C4" , x"CA" , x"5E" , x"5C" , x"A8" , x"E1" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5D" , x"D4" , x"BB" , x"5C" , x"60" , x"97" , x"E2" , x"8E" , x"E7" , x"8A" , x"5E" , x"66" , x"84" , x"F8" , x"F2" , x"F4" , x"F1" , x"FC" , x"B8" , x"DA" , x"B4" , x"5D" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5D" , x"AB" , x"DE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"76" , x"F1" , x"85" , x"66" , x"5E" , x"A3" , x"E4" , x"67" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7C" , x"F2" , x"7E" , x"66" , x"66" , x"5D" , x"DB" , x"B4" , x"9A" , x"EE" , x"80" , x"61" , x"66" , x"66" , x"61" , x"8A" , x"84" , x"80" , x"9C" , x"F3" , x"D9" , x"68" , x"57" , x"BE" , x"D1" , x"5D" , x"62" , x"99" , x"EC" , x"6C" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"63" , x"E2" , x"AB" , x"5D" , x"5E" , x"9F" , x"E0" , x"8D" , x"E7" , x"8A" , x"5E" , x"66" , x"83" , x"F8" , x"F7" , x"F8" , x"FA" , x"F4" , x"9A" , x"D5" , x"D8" , x"60" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5D" , x"AB" , x"DE" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"85" , x"66" , x"5E" , x"A3" , x"E4" , x"67" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F2" , x"7E" , x"66" , x"66" , x"5D" , x"DB" , x"B3" , x"8D" , x"F6" , x"AD" , x"5C" , x"66" , x"66" , x"6F" , x"CE" , x"C8" , x"BD" , x"E6" , x"FA" , x"A5" , x"5E" , x"5A" , x"B3" , x"DB" , x"5F" , x"66" , x"88" , x"F3" , x"7B" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"6F" , x"EE" , x"9A" , x"60" , x"5D" , x"AC" , x"DA" , x"8A" , x"E8" , x"8A" , x"5E" , x"66" , x"80" , x"EF" , x"B9" , x"B4" , x"B8" , x"AA" , x"79" , x"B0" , x"F1" , x"75" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"5D" , x"AB" , x"DE" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"85" , x"66" , x"5E" , x"A3" , x"E3" , x"67" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F3" , x"7E" , x"66" , x"66" , x"5D" , x"DB" , x"B2" , x"6F" , x"DB" , x"D9" , x"62" , x"65" , x"66" , x"60" , x"D6" , x"FD" , x"F8" , x"FE" , x"CA" , x"71" , x"63" , x"5C" , x"A2" , x"E5" , x"66" , x"66" , x"76" , x"F3" , x"90" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"66" , x"61" , x"82" , x"F4" , x"84" , x"66" , x"5D" , x"BE" , x"D0" , x"87" , x"E8" , x"89" , x"5E" , x"66" , x"7D" , x"EA" , x"8E" , x"7A" , x"7F" , x"73" , x"62" , x"88" , x"F5" , x"A2" , x"5B" , x"66" , x"65" , x"66" , x"66" , x"5D" , x"AB" , x"DE" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"74" , x"F1" , x"84" , x"66" , x"5E" , x"A3" , x"E3" , x"67" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F3" , x"7F" , x"66" , x"66" , x"5E" , x"DC" , x"B0" , x"57" , x"B0" , x"F4" , x"83" , x"5C" , x"66" , x"58" , x"A0" , x"F5" , x"F0" , x"CE" , x"8E" , x"5E" , x"66" , x"5B" , x"93" , x"ED" , x"6D" , x"66" , x"67" , x"E8" , x"B6" , x"5D" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5C" , x"A4" , x"F1" , x"70" , x"66" , x"5E" , x"CE" , x"C5" , x"82" , x"E9" , x"89" , x"5E" , x"66" , x"7D" , x"EF" , x"86" , x"5F" , x"62" , x"65" , x"66" , x"6C" , x"E2" , x"CE" , x"60" , x"66" , x"67" , x"66" , x"66" , x"5D" , x"AB" , x"DE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"84" , x"66" , x"5E" , x"A3" , x"E3" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F3" , x"7F" , x"66" , x"66" , x"5F" , x"DC" , x"B0" , x"55" , x"84" , x"F4" , x"B4" , x"5A" , x"66" , x"5C" , x"71" , x"E9" , x"CA" , x"89" , x"6A" , x"63" , x"67" , x"5F" , x"85" , x"F2" , x"78" , x"66" , x"5A" , x"D0" , x"DB" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5E" , x"CD" , x"DE" , x"62" , x"66" , x"62" , x"DF" , x"B4" , x"7A" , x"EA" , x"89" , x"5E" , x"66" , x"7C" , x"F2" , x"7D" , x"66" , x"66" , x"66" , x"67" , x"60" , x"BE" , x"EE" , x"72" , x"63" , x"66" , x"66" , x"66" , x"5D" , x"AB" , x"DE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"84" , x"66" , x"5E" , x"A3" , x"E3" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F3" , x"7E" , x"66" , x"66" , x"5F" , x"DC" , x"B1" , x"5B" , x"68" , x"DA" , x"DD" , x"68" , x"62" , x"65" , x"58" , x"CA" , x"E4" , x"85" , x"65" , x"66" , x"67" , x"65" , x"74" , x"F1" , x"8B" , x"62" , x"58" , x"AA" , x"F3" , x"89" , x"5C" , x"66" , x"66" , x"66" , x"5C" , x"7B" , x"EE" , x"BA" , x"5C" , x"66" , x"6A" , x"EB" , x"9D" , x"72" , x"EA" , x"89" , x"5E" , x"66" , x"7C" , x"F2" , x"7C" , x"66" , x"66" , x"66" , x"66" , x"60" , x"8D" , x"F7" , x"97" , x"5D" , x"66" , x"66" , x"66" , x"5D" , x"AB" , x"DE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"85" , x"66" , x"5D" , x"A3" , x"E3" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F3" , x"80" , x"66" , x"66" , x"60" , x"DB" , x"B2" , x"5D" , x"5E" , x"AE" , x"F6" , x"8D" , x"5C" , x"66" , x"57" , x"9B" , x"F8" , x"9D" , x"62" , x"66" , x"67" , x"66" , x"67" , x"E9" , x"A7" , x"5C" , x"5E" , x"7F" , x"F4" , x"BC" , x"67" , x"5B" , x"5E" , x"5A" , x"61" , x"AF" , x"FA" , x"8C" , x"60" , x"64" , x"79" , x"F2" , x"86" , x"6C" , x"EB" , x"88" , x"5F" , x"66" , x"7C" , x"F2" , x"7B" , x"66" , x"66" , x"66" , x"67" , x"65" , x"6C" , x"E8" , x"C5" , x"60" , x"66" , x"67" , x"66" , x"5D" , x"AB" , x"DE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"86" , x"66" , x"5D" , x"A3" , x"E3" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7E" , x"F3" , x"7F" , x"66" , x"66" , x"60" , x"DB" , x"B0" , x"5D" , x"63" , x"7C" , x"F2" , x"BC" , x"5A" , x"66" , x"60" , x"70" , x"E9" , x"CB" , x"63" , x"66" , x"67" , x"66" , x"5D" , x"D7" , x"C6" , x"5D" , x"66" , x"61" , x"D4" , x"F0" , x"91" , x"6C" , x"62" , x"6B" , x"88" , x"E7" , x"E3" , x"6D" , x"66" , x"5D" , x"96" , x"F2" , x"73" , x"70" , x"EF" , x"8A" , x"5F" , x"66" , x"7C" , x"F2" , x"7C" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"C6" , x"EA" , x"6F" , x"66" , x"67" , x"66" , x"5C" , x"AC" , x"DE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"85" , x"66" , x"5E" , x"A3" , x"E3" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7E" , x"F3" , x"7F" , x"66" , x"66" , x"60" , x"DC" , x"B0" , x"5C" , x"66" , x"61" , x"D4" , x"E3" , x"67" , x"62" , x"66" , x"5F" , x"C5" , x"EC" , x"76" , x"62" , x"67" , x"66" , x"57" , x"BF" , x"E0" , x"65" , x"66" , x"59" , x"A1" , x"FB" , x"D9" , x"95" , x"86" , x"91" , x"CF" , x"FD" , x"AF" , x"5F" , x"66" , x"5A" , x"BA" , x"E7" , x"64" , x"74" , x"F0" , x"89" , x"5F" , x"66" , x"7D" , x"F2" , x"7B" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5E" , x"99" , x"F7" , x"8D" , x"61" , x"66" , x"66" , x"5C" , x"AC" , x"DE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"85" , x"66" , x"5E" , x"A3" , x"E3" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7C" , x"F3" , x"80" , x"66" , x"66" , x"5F" , x"DC" , x"AF" , x"5C" , x"66" , x"5C" , x"A5" , x"F7" , x"8F" , x"5A" , x"66" , x"5C" , x"94" , x"F8" , x"A2" , x"5D" , x"66" , x"66" , x"58" , x"9E" , x"F0" , x"76" , x"64" , x"60" , x"6E" , x"D0" , x"FE" , x"E8" , x"D5" , x"E4" , x"FE" , x"DB" , x"77" , x"61" , x"66" , x"60" , x"D8" , x"CE" , x"5B" , x"75" , x"F0" , x"8A" , x"5F" , x"66" , x"7D" , x"F2" , x"7B" , x"66" , x"66" , x"66" , x"66" , x"66" , x"63" , x"73" , x"ED" , x"BD" , x"62" , x"66" , x"66" , x"5C" , x"AD" , x"DE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"74" , x"F1" , x"85" , x"66" , x"5D" , x"A3" , x"E3" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F3" , x"80" , x"66" , x"66" , x"60" , x"DB" , x"AF" , x"5D" , x"66" , x"60" , x"78" , x"EF" , x"C0" , x"5A" , x"66" , x"62" , x"6A" , x"E7" , x"CE" , x"5E" , x"66" , x"66" , x"5B" , x"79" , x"F3" , x"9F" , x"5D" , x"66" , x"5C" , x"93" , x"E2" , x"FD" , x"FC" , x"FE" , x"E8" , x"9C" , x"5E" , x"66" , x"5F" , x"74" , x"ED" , x"AB" , x"59" , x"76" , x"EF" , x"89" , x"60" , x"66" , x"7D" , x"F2" , x"7B" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"62" , x"CF" , x"E4" , x"6D" , x"66" , x"66" , x"5B" , x"AD" , x"DE" , x"62" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"85" , x"66" , x"5D" , x"A3" , x"E3" , x"65" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F3" , x"7E" , x"66" , x"66" , x"60" , x"DC" , x"AF" , x"5D" , x"66" , x"66" , x"61" , x"CE" , x"E5" , x"6E" , x"61" , x"66" , x"60" , x"C2" , x"EE" , x"74" , x"5E" , x"66" , x"65" , x"64" , x"E3" , x"C9" , x"60" , x"66" , x"60" , x"65" , x"95" , x"C7" , x"DF" , x"CD" , x"9C" , x"6A" , x"5F" , x"66" , x"56" , x"9E" , x"F3" , x"83" , x"5D" , x"75" , x"EF" , x"89" , x"60" , x"66" , x"7C" , x"F2" , x"7B" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"5E" , x"A3" , x"F5" , x"86" , x"61" , x"66" , x"5A" , x"AD" , x"DE" , x"62" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"74" , x"F1" , x"85" , x"66" , x"5D" , x"A3" , x"E3" , x"65" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F3" , x"7F" , x"66" , x"66" , x"60" , x"DB" , x"AF" , x"5D" , x"66" , x"66" , x"5C" , x"9D" , x"F7" , x"99" , x"5C" , x"66" , x"5F" , x"92" , x"F7" , x"A4" , x"5A" , x"66" , x"66" , x"5A" , x"C4" , x"E9" , x"74" , x"60" , x"66" , x"57" , x"6F" , x"82" , x"8C" , x"85" , x"74" , x"57" , x"66" , x"63" , x"5B" , x"CA" , x"E7" , x"69" , x"66" , x"73" , x"EE" , x"8A" , x"61" , x"66" , x"7B" , x"F1" , x"7C" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"63" , x"78" , x"F0" , x"B4" , x"5F" , x"66" , x"5B" , x"AD" , x"DE" , x"62" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"86" , x"66" , x"5D" , x"A3" , x"E3" , x"65" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F3" , x"7F" , x"66" , x"66" , x"60" , x"DB" , x"AE" , x"5C" , x"66" , x"67" , x"62" , x"72" , x"EB" , x"C6" , x"5D" , x"66" , x"64" , x"6B" , x"E4" , x"D3" , x"61" , x"66" , x"66" , x"59" , x"98" , x"F8" , x"A3" , x"5C" , x"66" , x"66" , x"56" , x"5A" , x"68" , x"5C" , x"51" , x"63" , x"66" , x"58" , x"80" , x"ED" , x"C4" , x"5D" , x"66" , x"70" , x"EE" , x"8B" , x"60" , x"66" , x"7C" , x"F1" , x"7C" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"65" , x"D7" , x"DC" , x"66" , x"66" , x"5B" , x"AD" , x"DE" , x"62" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"85" , x"66" , x"5D" , x"A4" , x"E3" , x"65" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F3" , x"7F" , x"66" , x"66" , x"61" , x"DB" , x"AF" , x"5C" , x"66" , x"67" , x"66" , x"62" , x"CA" , x"E9" , x"6F" , x"60" , x"66" , x"5E" , x"BB" , x"F0" , x"7B" , x"5D" , x"66" , x"5F" , x"6E" , x"E7" , x"D1" , x"68" , x"60" , x"66" , x"66" , x"5C" , x"55" , x"59" , x"66" , x"66" , x"62" , x"58" , x"AD" , x"F8" , x"93" , x"5C" , x"66" , x"71" , x"EE" , x"89" , x"60" , x"66" , x"7C" , x"F1" , x"7D" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"AD" , x"F2" , x"7F" , x"64" , x"5C" , x"AE" , x"DE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"F1" , x"84" , x"66" , x"5D" , x"A4" , x"E2" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F3" , x"7E" , x"66" , x"66" , x"61" , x"DB" , x"AF" , x"5C" , x"66" , x"66" , x"66" , x"61" , x"9B" , x"F8" , x"9C" , x"5A" , x"66" , x"5F" , x"88" , x"F6" , x"AA" , x"58" , x"66" , x"66" , x"5B" , x"BE" , x"F7" , x"97" , x"5C" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"58" , x"7E" , x"E2" , x"E1" , x"6B" , x"62" , x"66" , x"71" , x"EE" , x"8A" , x"5E" , x"66" , x"7C" , x"F1" , x"7D" , x"66" , x"67" , x"66" , x"66" , x"66" , x"67" , x"66" , x"62" , x"81" , x"F3" , x"AC" , x"5F" , x"5C" , x"AF" , x"DE" , x"62" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"74" , x"F2" , x"84" , x"66" , x"5D" , x"A4" , x"E2" , x"65" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F2" , x"7E" , x"66" , x"66" , x"62" , x"DC" , x"AF" , x"5D" , x"66" , x"66" , x"66" , x"64" , x"71" , x"E8" , x"CB" , x"5D" , x"66" , x"66" , x"6D" , x"E1" , x"D5" , x"5E" , x"62" , x"66" , x"5A" , x"8B" , x"F4" , x"D0" , x"79" , x"5D" , x"5F" , x"66" , x"66" , x"66" , x"60" , x"57" , x"68" , x"B0" , x"FD" , x"AF" , x"5B" , x"66" , x"66" , x"72" , x"EE" , x"89" , x"5F" , x"66" , x"7C" , x"F1" , x"7E" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"69" , x"DE" , x"D5" , x"63" , x"5B" , x"B0" , x"DE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"ED" , x"85" , x"62" , x"5D" , x"A7" , x"E0" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"F0" , x"82" , x"58" , x"5C" , x"61" , x"DB" , x"AF" , x"5C" , x"66" , x"66" , x"67" , x"66" , x"61" , x"C3" , x"EE" , x"78" , x"5B" , x"66" , x"65" , x"BB" , x"F3" , x"81" , x"5A" , x"66" , x"62" , x"63" , x"C7" , x"FC" , x"AB" , x"75" , x"57" , x"4A" , x"4B" , x"48" , x"4E" , x"6D" , x"92" , x"ED" , x"E5" , x"7C" , x"5D" , x"66" , x"66" , x"72" , x"ED" , x"8B" , x"5B" , x"5E" , x"7C" , x"EF" , x"7D" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"B6" , x"EF" , x"79" , x"53" , x"B0" , x"DE" , x"62" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"75" , x"EC" , x"90" , x"64" , x"64" , x"B3" , x"DC" , x"64" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7D" , x"ED" , x"8E" , x"6E" , x"6F" , x"76" , x"D8" , x"AE" , x"5D" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"91" , x"F7" , x"A2" , x"60" , x"64" , x"71" , x"9A" , x"F3" , x"AF" , x"57" , x"66" , x"66" , x"5A" , x"90" , x"ED" , x"F0" , x"A1" , x"7A" , x"71" , x"70" , x"6F" , x"76" , x"90" , x"DB" , x"FC" , x"AF" , x"5E" , x"65" , x"67" , x"66" , x"73" , x"EB" , x"96" , x"61" , x"61" , x"89" , x"EC" , x"7D" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"88" , x"F6" , x"9F" , x"61" , x"B3" , x"DE" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"70" , x"EB" , x"9D" , x"81" , x"7E" , x"C4" , x"D1" , x"61" , x"66" , x"66" , x"66" , x"67" , x"66" , x"7C" , x"EC" , x"96" , x"8B" , x"8F" , x"87" , x"D7" , x"AD" , x"5D" , x"66" , x"66" , x"66" , x"66" , x"64" , x"6B" , x"E5" , x"CC" , x"7E" , x"86" , x"87" , x"86" , x"D4" , x"DB" , x"5D" , x"66" , x"66" , x"61" , x"64" , x"B4" , x"FB" , x"ED" , x"B5" , x"91" , x"8D" , x"8F" , x"A5" , x"DE" , x"FE" , x"D1" , x"77" , x"60" , x"66" , x"67" , x"66" , x"72" , x"E9" , x"9C" , x"7F" , x"81" , x"91" , x"EB" , x"7D" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"6A" , x"E5" , x"C9" , x"75" , x"B4" , x"DD" , x"62" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"E3" , x"DB" , x"CB" , x"C9" , x"EC" , x"B9" , x"5F" , x"66" , x"66" , x"66" , x"67" , x"66" , x"76" , x"EF" , x"DF" , x"DB" , x"DD" , x"D8" , x"F4" , x"A3" , x"5E" , x"66" , x"66" , x"66" , x"67" , x"66" , x"5E" , x"BC" , x"F2" , x"C7" , x"CA" , x"CC" , x"C8" , x"E0" , x"E5" , x"66" , x"66" , x"67" , x"66" , x"5C" , x"7E" , x"C9" , x"FE" , x"F7" , x"E4" , x"DB" , x"E0" , x"F3" , x"FF" , x"E0" , x"92" , x"60" , x"66" , x"66" , x"67" , x"66" , x"6C" , x"E7" , x"D9" , x"CB" , x"CC" , x"D4" , x"F0" , x"77" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"BF" , x"F0" , x"C6" , x"E5" , x"D2" , x"60" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"CD" , x"FD" , x"FB" , x"FA" , x"FC" , x"99" , x"60" , x"66" , x"67" , x"66" , x"66" , x"66" , x"69" , x"E1" , x"FD" , x"FC" , x"FD" , x"FE" , x"FC" , x"8A" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5E" , x"8A" , x"F2" , x"FD" , x"FD" , x"FC" , x"FA" , x"FD" , x"E4" , x"69" , x"66" , x"66" , x"66" , x"65" , x"5E" , x"88" , x"C6" , x"F5" , x"FC" , x"FD" , x"FD" , x"F9" , x"D9" , x"97" , x"69" , x"64" , x"66" , x"66" , x"66" , x"66" , x"62" , x"D5" , x"FD" , x"FB" , x"FB" , x"FD" , x"E2" , x"69" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"92" , x"F5" , x"FB" , x"FE" , x"B7" , x"5D" , x"66" , x"65" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5E" , x"9E" , x"E5" , x"E3" , x"E7" , x"D6" , x"79" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"63" , x"AD" , x"DC" , x"D7" , x"D7" , x"DD" , x"C9" , x"6F" , x"66" , x"67" , x"66" , x"66" , x"66" , x"67" , x"64" , x"6B" , x"D6" , x"EA" , x"E6" , x"E6" , x"E4" , x"EB" , x"D8" , x"69" , x"66" , x"66" , x"66" , x"66" , x"61" , x"63" , x"85" , x"A8" , x"CF" , x"D9" , x"D4" , x"B6" , x"8C" , x"6C" , x"60" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"A3" , x"E7" , x"E3" , x"E3" , x"E7" , x"AF" , x"62" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"64" , x"71" , x"D9" , x"E8" , x"DF" , x"87" , x"60" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"63" , x"6E" , x"95" , x"94" , x"95" , x"8E" , x"69" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"64" , x"76" , x"8D" , x"89" , x"8A" , x"8C" , x"85" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"63" , x"96" , x"97" , x"92" , x"93" , x"94" , x"96" , x"91" , x"65" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"5E" , x"77" , x"85" , x"8B" , x"88" , x"7E" , x"66" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"65" , x"66" , x"62" , x"71" , x"94" , x"93" , x"93" , x"95" , x"75" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"94" , x"95" , x"93" , x"6A" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"60" , x"6A" , x"72" , x"70" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"63" , x"67" , x"65" , x"63" , x"67" , x"65" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"65" , x"66" , x"63" , x"67" , x"79" , x"76" , x"75" , x"73" , x"75" , x"66" , x"65" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"62" , x"5A" , x"5F" , x"62" , x"63" , x"5E" , x"61" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5D" , x"70" , x"76" , x"75" , x"6D" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"65" , x"66" , x"65" , x"66" , x"77" , x"68" , x"64" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5E" , x"5C" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"63" , x"61" , x"62" , x"63" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5F" , x"55" , x"55" , x"5A" , x"5B" , x"5B" , x"62" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"62" , x"5F" , x"61" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"5A" , x"57" , x"58" , x"5E" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"62" , x"58" , x"5F" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"66" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"67" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"65" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ),
( x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" , x"66" ) 
);

CONSTANT Plantilla_TronB : ImageMatrix(0 TO 99, 0 TO 99) := (
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"FE" , x"FF" , x"FF" , x"FE" , x"FD" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"FE" , x"FF" , x"FE" , x"FD" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FD" , x"FB" , x"FB" , x"FD" , x"FD" , x"FE" , x"FD" , x"FD" , x"FE" , x"FD" , x"FE" , x"FE" , x"FE" , x"FD" , x"FB" , x"F9" , x"F8" , x"FB" , x"FD" , x"FA" , x"FA" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"F9" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"B8" , x"8E" , x"89" , x"8A" , x"8D" , x"93" , x"9A" , x"B2" , x"F3" , x"FF" , x"FF" , x"FA" , x"C2" , x"9F" , x"8C" , x"89" , x"89" , x"87" , x"87" , x"86" , x"8A" , x"8B" , x"8A" , x"8B" , x"8B" , x"8B" , x"8A" , x"8B" , x"8B" , x"89" , x"88" , x"86" , x"84" , x"87" , x"89" , x"86" , x"85" , x"8C" , x"A4" , x"CE" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FE" , x"CA" , x"A3" , x"90" , x"94" , x"B7" , x"EF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"E4" , x"A3" , x"8A" , x"B7" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"F7" , x"A5" , x"8A" , x"84" , x"8C" , x"9E" , x"E9" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FD" , x"FF" , x"C6" , x"7E" , x"8F" , x"8E" , x"8F" , x"8F" , x"8F" , x"8E" , x"90" , x"A3" , x"FF" , x"F9" , x"95" , x"86" , x"8D" , x"8D" , x"8E" , x"8E" , x"8E" , x"8E" , x"8F" , x"8F" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8E" , x"8F" , x"8C" , x"7C" , x"A3" , x"FA" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"EE" , x"93" , x"78" , x"88" , x"8D" , x"89" , x"81" , x"83" , x"D8" , x"FF" , x"FE" , x"FF" , x"FF" , x"FE" , x"FF" , x"FA" , x"88" , x"90" , x"8F" , x"84" , x"D3" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FF" , x"B5" , x"80" , x"8F" , x"8D" , x"8E" , x"8F" , x"8F" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FE" , x"FF" , x"99" , x"B9" , x"DD" , x"D5" , x"D8" , x"D8" , x"D6" , x"DA" , x"D1" , x"83" , x"F8" , x"BA" , x"89" , x"BE" , x"D5" , x"D6" , x"D6" , x"D6" , x"D6" , x"D7" , x"D8" , x"D7" , x"D7" , x"D6" , x"D6" , x"D7" , x"D6" , x"D6" , x"D7" , x"D7" , x"D6" , x"D6" , x"D6" , x"D6" , x"D6" , x"D6" , x"D6" , x"D7" , x"D9" , x"D1" , x"AD" , x"89" , x"A1" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"F5" , x"85" , x"8A" , x"A8" , x"CD" , x"D7" , x"D3" , x"B7" , x"92" , x"7A" , x"DA" , x"FF" , x"FE" , x"FF" , x"FD" , x"FF" , x"D9" , x"93" , x"D5" , x"DE" , x"C5" , x"9D" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"90" , x"BB" , x"DC" , x"D4" , x"D7" , x"D3" , x"86" , x"E1" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"92" , x"EF" , x"FF" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"A1" , x"D1" , x"8E" , x"C4" , x"FF" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"F5" , x"C1" , x"7A" , x"D0" , x"FF" , x"FD" , x"FF" , x"FF" , x"FE" , x"FF" , x"9A" , x"8C" , x"C6" , x"F4" , x"FD" , x"FF" , x"FF" , x"FA" , x"D7" , x"9A" , x"7D" , x"F2" , x"FE" , x"FE" , x"FD" , x"FF" , x"BF" , x"CA" , x"FF" , x"FF" , x"F2" , x"8E" , x"F6" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FE" , x"91" , x"F1" , x"FF" , x"FF" , x"FD" , x"FF" , x"B5" , x"C5" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"FB" , x"98" , x"F6" , x"EB" , x"EB" , x"EA" , x"EA" , x"EB" , x"E6" , x"F8" , x"BA" , x"8E" , x"9B" , x"F6" , x"F8" , x"E7" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"EA" , x"E9" , x"EF" , x"FC" , x"FA" , x"AF" , x"8F" , x"FF" , x"FE" , x"FF" , x"FD" , x"FF" , x"CF" , x"7F" , x"C9" , x"FF" , x"FD" , x"F0" , x"E8" , x"ED" , x"FA" , x"FF" , x"DF" , x"92" , x"A5" , x"FF" , x"FD" , x"FD" , x"FF" , x"B6" , x"E6" , x"F4" , x"E7" , x"F9" , x"A5" , x"D5" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F7" , x"9F" , x"FB" , x"EB" , x"EA" , x"E8" , x"F7" , x"D4" , x"BD" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F6" , x"9A" , x"EE" , x"A1" , x"99" , x"98" , x"99" , x"9B" , x"93" , x"D3" , x"C5" , x"67" , x"C1" , x"FE" , x"B8" , x"97" , x"99" , x"97" , x"97" , x"97" , x"97" , x"99" , x"99" , x"99" , x"99" , x"99" , x"9A" , x"9B" , x"9A" , x"99" , x"9A" , x"9B" , x"99" , x"99" , x"98" , x"97" , x"98" , x"99" , x"99" , x"99" , x"A0" , x"C6" , x"FD" , x"E7" , x"85" , x"E2" , x"FF" , x"FD" , x"FF" , x"F9" , x"84" , x"B6" , x"FB" , x"F6" , x"C9" , x"A2" , x"9E" , x"A1" , x"BB" , x"EC" , x"FF" , x"CF" , x"7C" , x"E4" , x"FE" , x"FC" , x"FF" , x"AF" , x"EC" , x"B3" , x"94" , x"E8" , x"D4" , x"B2" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F4" , x"A9" , x"EB" , x"9A" , x"9F" , x"96" , x"C2" , x"DC" , x"BA" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F5" , x"98" , x"F0" , x"8F" , x"71" , x"73" , x"79" , x"87" , x"81" , x"D0" , x"CA" , x"82" , x"E9" , x"D8" , x"81" , x"74" , x"72" , x"71" , x"72" , x"72" , x"72" , x"72" , x"73" , x"73" , x"72" , x"72" , x"72" , x"73" , x"72" , x"72" , x"73" , x"73" , x"72" , x"72" , x"71" , x"70" , x"71" , x"72" , x"72" , x"73" , x"78" , x"88" , x"C4" , x"FF" , x"B8" , x"B3" , x"FF" , x"FB" , x"FF" , x"BE" , x"93" , x"EE" , x"F9" , x"B3" , x"88" , x"7A" , x"73" , x"78" , x"85" , x"9F" , x"E9" , x"FF" , x"B0" , x"A1" , x"FF" , x"FD" , x"FF" , x"A8" , x"F1" , x"A7" , x"82" , x"C5" , x"F3" , x"99" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F2" , x"AA" , x"EA" , x"85" , x"8E" , x"7D" , x"BA" , x"DF" , x"BA" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F4" , x"9A" , x"F5" , x"9A" , x"D9" , x"DE" , x"E4" , x"F5" , x"C2" , x"D1" , x"CA" , x"9C" , x"F7" , x"A5" , x"9B" , x"C9" , x"D2" , x"CD" , x"CC" , x"C8" , x"C8" , x"C3" , x"BB" , x"BA" , x"BE" , x"C5" , x"C7" , x"C6" , x"C4" , x"C0" , x"BC" , x"BF" , x"C8" , x"D0" , x"D4" , x"D4" , x"D1" , x"CE" , x"CB" , x"C6" , x"C1" , x"94" , x"88" , x"E8" , x"E6" , x"94" , x"FF" , x"FF" , x"F9" , x"7F" , x"C7" , x"FF" , x"BE" , x"7F" , x"91" , x"B6" , x"BC" , x"B5" , x"99" , x"73" , x"A2" , x"F7" , x"E5" , x"84" , x"EA" , x"FF" , x"FF" , x"A2" , x"F5" , x"AE" , x"D0" , x"A0" , x"FC" , x"9E" , x"E2" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F0" , x"AB" , x"EF" , x"9B" , x"F9" , x"C0" , x"B9" , x"E3" , x"BA" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F3" , x"9A" , x"F7" , x"AB" , x"FF" , x"FF" , x"FF" , x"FF" , x"D5" , x"CE" , x"C8" , x"B4" , x"F0" , x"95" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"92" , x"B7" , x"F9" , x"90" , x"E9" , x"FF" , x"C8" , x"8F" , x"F6" , x"DF" , x"86" , x"AB" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"C7" , x"79" , x"C0" , x"FF" , x"B3" , x"B4" , x"FF" , x"FF" , x"9D" , x"F5" , x"A7" , x"FF" , x"9D" , x"F0" , x"C9" , x"B6" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F0" , x"AA" , x"EF" , x"A9" , x"FF" , x"DA" , x"B3" , x"E3" , x"BB" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F3" , x"9A" , x"F7" , x"AA" , x"FD" , x"FD" , x"FC" , x"FE" , x"D0" , x"CE" , x"C6" , x"C8" , x"E0" , x"B2" , x"FF" , x"FB" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FB" , x"FF" , x"E0" , x"8A" , x"F4" , x"AD" , x"CA" , x"FF" , x"8F" , x"C1" , x"FF" , x"A9" , x"93" , x"FF" , x"FD" , x"FB" , x"FD" , x"FC" , x"FB" , x"FF" , x"B0" , x"8D" , x"EE" , x"E3" , x"8D" , x"FB" , x"FF" , x"9A" , x"F4" , x"A3" , x"FF" , x"B1" , x"CF" , x"EA" , x"93" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F0" , x"AC" , x"EF" , x"A8" , x"FE" , x"D9" , x"B2" , x"E5" , x"BC" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F3" , x"9B" , x"F7" , x"AD" , x"FE" , x"FC" , x"FB" , x"FD" , x"D1" , x"CE" , x"C6" , x"D5" , x"C7" , x"CA" , x"FE" , x"FD" , x"FE" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FE" , x"FE" , x"FE" , x"FE" , x"FD" , x"FE" , x"FE" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"99" , x"E2" , x"CC" , x"B3" , x"F6" , x"76" , x"EA" , x"DF" , x"83" , x"EA" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FC" , x"FB" , x"82" , x"BC" , x"FF" , x"93" , x"D9" , x"FF" , x"94" , x"F4" , x"A2" , x"FF" , x"D4" , x"A3" , x"FB" , x"94" , x"DE" , x"FF" , x"FE" , x"FF" , x"FF" , x"FE" , x"FF" , x"F1" , x"AB" , x"EF" , x"A8" , x"FF" , x"DA" , x"B3" , x"E5" , x"BD" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F3" , x"9B" , x"F7" , x"A7" , x"FF" , x"FF" , x"FF" , x"FF" , x"D9" , x"CF" , x"C8" , x"DC" , x"AC" , x"DD" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"C6" , x"CB" , x"DF" , x"A9" , x"CC" , x"99" , x"FF" , x"B0" , x"AF" , x"FF" , x"FF" , x"E1" , x"9B" , x"85" , x"99" , x"E0" , x"FF" , x"FF" , x"CA" , x"8B" , x"F7" , x"C4" , x"AC" , x"FF" , x"92" , x"F4" , x"A4" , x"F9" , x"F7" , x"8D" , x"F5" , x"C1" , x"B2" , x"FF" , x"FD" , x"FF" , x"FF" , x"FE" , x"FF" , x"F2" , x"AB" , x"EF" , x"A7" , x"FF" , x"DA" , x"B3" , x"E5" , x"BF" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F3" , x"98" , x"F2" , x"8F" , x"98" , x"9F" , x"A5" , x"B3" , x"9A" , x"D2" , x"CB" , x"E2" , x"A1" , x"E6" , x"FF" , x"FF" , x"E6" , x"AE" , x"A5" , x"9E" , x"9D" , x"9E" , x"9B" , x"94" , x"93" , x"9B" , x"A3" , x"A0" , x"97" , x"95" , x"92" , x"90" , x"90" , x"93" , x"96" , x"95" , x"8A" , x"86" , x"8A" , x"8C" , x"8E" , x"97" , x"B1" , x"9C" , x"B9" , x"EB" , x"A5" , x"A8" , x"C8" , x"F2" , x"88" , x"EA" , x"FF" , x"D6" , x"74" , x"84" , x"88" , x"86" , x"78" , x"D7" , x"FF" , x"FD" , x"88" , x"D5" , x"E9" , x"91" , x"FF" , x"96" , x"F4" , x"A3" , x"F2" , x"FF" , x"A1" , x"D9" , x"E6" , x"92" , x"FF" , x"FE" , x"FF" , x"FF" , x"FE" , x"FF" , x"F2" , x"AB" , x"EF" , x"A5" , x"FF" , x"DA" , x"B1" , x"E5" , x"BF" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F4" , x"9A" , x"EE" , x"91" , x"82" , x"84" , x"84" , x"83" , x"83" , x"CD" , x"CD" , x"E4" , x"9B" , x"EA" , x"FF" , x"F7" , x"7F" , x"83" , x"85" , x"85" , x"85" , x"85" , x"85" , x"85" , x"85" , x"85" , x"85" , x"85" , x"85" , x"85" , x"85" , x"85" , x"85" , x"85" , x"85" , x"84" , x"85" , x"84" , x"84" , x"85" , x"85" , x"85" , x"84" , x"84" , x"AB" , x"EE" , x"88" , x"81" , x"E5" , x"D4" , x"9D" , x"FF" , x"E8" , x"75" , x"91" , x"B7" , x"CB" , x"BC" , x"95" , x"7B" , x"ED" , x"FE" , x"BF" , x"AB" , x"F7" , x"8D" , x"EC" , x"9E" , x"F5" , x"A4" , x"F3" , x"FF" , x"CC" , x"AB" , x"FA" , x"8C" , x"E3" , x"FF" , x"FE" , x"FF" , x"FE" , x"FF" , x"F2" , x"AB" , x"EF" , x"A3" , x"FF" , x"D9" , x"B1" , x"E5" , x"C0" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"F6" , x"96" , x"F1" , x"BE" , x"BC" , x"BD" , x"BC" , x"BD" , x"B6" , x"DE" , x"CC" , x"E5" , x"99" , x"EA" , x"FF" , x"C5" , x"89" , x"BC" , x"BD" , x"BC" , x"BD" , x"BD" , x"BD" , x"BD" , x"BC" , x"BC" , x"BC" , x"BC" , x"BC" , x"BC" , x"BD" , x"BD" , x"BC" , x"BC" , x"BC" , x"BC" , x"BC" , x"BC" , x"BC" , x"BC" , x"BC" , x"BC" , x"BD" , x"B9" , x"C6" , x"EC" , x"6C" , x"7B" , x"F5" , x"A9" , x"CE" , x"FF" , x"95" , x"8C" , x"D5" , x"FC" , x"FE" , x"FD" , x"DC" , x"94" , x"A3" , x"FF" , x"EF" , x"8C" , x"F5" , x"AB" , x"CC" , x"A4" , x"F6" , x"A4" , x"F6" , x"FF" , x"F3" , x"91" , x"F7" , x"B6" , x"B7" , x"FF" , x"FD" , x"FF" , x"FE" , x"FF" , x"F2" , x"AD" , x"EF" , x"A0" , x"FF" , x"DA" , x"B1" , x"E4" , x"C0" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FE" , x"FF" , x"FC" , x"91" , x"F7" , x"FD" , x"FB" , x"FB" , x"FB" , x"FB" , x"FA" , x"FE" , x"BF" , x"E7" , x"98" , x"ED" , x"FF" , x"99" , x"C1" , x"FF" , x"F9" , x"FB" , x"FB" , x"FB" , x"FB" , x"FB" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FB" , x"FB" , x"FB" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FA" , x"FD" , x"EA" , x"77" , x"A0" , x"F8" , x"93" , x"FA" , x"EC" , x"70" , x"C4" , x"FF" , x"F8" , x"EE" , x"F7" , x"FF" , x"D1" , x"79" , x"E9" , x"FF" , x"9D" , x"E3" , x"CF" , x"B3" , x"A6" , x"F6" , x"A6" , x"F7" , x"FF" , x"FF" , x"A3" , x"E0" , x"DF" , x"95" , x"FF" , x"FE" , x"FF" , x"FE" , x"FF" , x"F2" , x"AB" , x"EF" , x"A2" , x"FF" , x"DA" , x"B1" , x"E4" , x"BF" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"91" , x"DE" , x"FF" , x"F8" , x"F8" , x"F8" , x"F9" , x"FB" , x"F1" , x"AA" , x"EB" , x"99" , x"F2" , x"FF" , x"8C" , x"EA" , x"FB" , x"F6" , x"F8" , x"F8" , x"F8" , x"F8" , x"F8" , x"F8" , x"F7" , x"F7" , x"F7" , x"F7" , x"F7" , x"F8" , x"F8" , x"F8" , x"F7" , x"F7" , x"F7" , x"F7" , x"F7" , x"F7" , x"F7" , x"F7" , x"F7" , x"F8" , x"F7" , x"FC" , x"E9" , x"7F" , x"C1" , x"EC" , x"A5" , x"FF" , x"B9" , x"99" , x"F8" , x"F0" , x"B8" , x"9C" , x"B2" , x"EC" , x"FF" , x"A5" , x"B8" , x"FE" , x"BF" , x"C3" , x"EA" , x"A0" , x"A6" , x"F6" , x"A6" , x"F7" , x"FF" , x"FE" , x"C8" , x"B7" , x"F8" , x"89" , x"E9" , x"FF" , x"FE" , x"FE" , x"FF" , x"F1" , x"AB" , x"EF" , x"A5" , x"FF" , x"DA" , x"B3" , x"E4" , x"C0" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FD" , x"FF" , x"AD" , x"9C" , x"B5" , x"B1" , x"B1" , x"B1" , x"B1" , x"B3" , x"A6" , x"9B" , x"EE" , x"9A" , x"F7" , x"F8" , x"94" , x"F8" , x"BF" , x"AE" , x"B2" , x"B1" , x"B1" , x"B1" , x"B1" , x"AF" , x"B0" , x"B0" , x"B0" , x"B1" , x"B2" , x"B1" , x"B0" , x"B2" , x"B0" , x"B0" , x"B0" , x"B0" , x"B0" , x"B0" , x"B0" , x"B0" , x"B0" , x"B0" , x"B0" , x"B2" , x"AB" , x"85" , x"D8" , x"D1" , x"C1" , x"FF" , x"96" , x"CF" , x"FF" , x"AC" , x"82" , x"74" , x"7E" , x"A0" , x"FA" , x"DC" , x"97" , x"FF" , x"E1" , x"A1" , x"F7" , x"8A" , x"8E" , x"F4" , x"A4" , x"F7" , x"FF" , x"FF" , x"EF" , x"93" , x"FB" , x"AF" , x"C3" , x"FF" , x"FD" , x"FE" , x"FF" , x"F0" , x"AA" , x"EF" , x"A9" , x"FF" , x"DA" , x"B3" , x"E4" , x"C0" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FE" , x"FF" , x"EA" , x"7B" , x"7F" , x"7C" , x"7D" , x"7C" , x"7A" , x"7C" , x"79" , x"95" , x"F1" , x"9A" , x"F9" , x"F0" , x"9E" , x"F0" , x"8B" , x"7B" , x"7E" , x"7E" , x"7D" , x"7D" , x"7F" , x"7F" , x"7E" , x"7E" , x"80" , x"7E" , x"81" , x"7D" , x"7A" , x"80" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7F" , x"7A" , x"80" , x"E9" , x"B0" , x"DC" , x"FD" , x"8B" , x"F5" , x"D4" , x"7A" , x"A6" , x"CC" , x"9E" , x"71" , x"C5" , x"FB" , x"94" , x"F4" , x"FC" , x"99" , x"F9" , x"89" , x"75" , x"F1" , x"A3" , x"F8" , x"FF" , x"FE" , x"FF" , x"9D" , x"E6" , x"D9" , x"A3" , x"FF" , x"FD" , x"FE" , x"FF" , x"EF" , x"AB" , x"EF" , x"AB" , x"FF" , x"DA" , x"B3" , x"E4" , x"C1" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"E5" , x"C6" , x"C4" , x"BF" , x"C5" , x"C6" , x"C2" , x"DD" , x"AB" , x"F6" , x"9D" , x"FB" , x"ED" , x"A5" , x"EB" , x"93" , x"B3" , x"B3" , x"BB" , x"BD" , x"BF" , x"AD" , x"6C" , x"64" , x"63" , x"6C" , x"CE" , x"ED" , x"E0" , x"DD" , x"9B" , x"63" , x"63" , x"62" , x"62" , x"61" , x"62" , x"62" , x"62" , x"61" , x"62" , x"61" , x"63" , x"5A" , x"80" , x"F3" , x"9E" , x"F7" , x"E0" , x"A0" , x"FB" , x"A1" , x"A9" , x"FF" , x"FF" , x"FF" , x"A8" , x"94" , x"F9" , x"B1" , x"D5" , x"FF" , x"A2" , x"F2" , x"A4" , x"7B" , x"F0" , x"A4" , x"F7" , x"FF" , x"FC" , x"FE" , x"BF" , x"BF" , x"F4" , x"93" , x"FA" , x"FF" , x"FE" , x"FD" , x"F1" , x"AD" , x"F0" , x"AF" , x"FF" , x"DA" , x"B3" , x"E4" , x"C0" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"AE" , x"F6" , x"9C" , x"FC" , x"EE" , x"AC" , x"EB" , x"BE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"9A" , x"76" , x"70" , x"74" , x"A1" , x"C5" , x"FF" , x"FF" , x"B6" , x"75" , x"71" , x"71" , x"71" , x"70" , x"72" , x"72" , x"71" , x"6F" , x"71" , x"71" , x"71" , x"69" , x"95" , x"F5" , x"9F" , x"FF" , x"C2" , x"CB" , x"EA" , x"86" , x"F5" , x"FF" , x"FC" , x"FF" , x"F9" , x"85" , x"DD" , x"D9" , x"B9" , x"FF" , x"B1" , x"E5" , x"BA" , x"83" , x"EF" , x"A3" , x"F6" , x"FF" , x"FD" , x"FF" , x"E4" , x"96" , x"FC" , x"A4" , x"DB" , x"FE" , x"FF" , x"FF" , x"FD" , x"AD" , x"F0" , x"B0" , x"FF" , x"DA" , x"B3" , x"E4" , x"C1" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FC" , x"FE" , x"AA" , x"F6" , x"9F" , x"FC" , x"EE" , x"AD" , x"EC" , x"C1" , x"FD" , x"FB" , x"FD" , x"FC" , x"FD" , x"E1" , x"88" , x"98" , x"95" , x"97" , x"9B" , x"97" , x"D6" , x"ED" , x"8B" , x"9B" , x"95" , x"94" , x"96" , x"98" , x"96" , x"95" , x"94" , x"93" , x"95" , x"95" , x"93" , x"8C" , x"AD" , x"EF" , x"A5" , x"FF" , x"A8" , x"E7" , x"CB" , x"AF" , x"FF" , x"FD" , x"FF" , x"FD" , x"FF" , x"B9" , x"B8" , x"F2" , x"AD" , x"FF" , x"C3" , x"D4" , x"CC" , x"8C" , x"EE" , x"A2" , x"F5" , x"FF" , x"FF" , x"FF" , x"FE" , x"96" , x"ED" , x"D0" , x"B4" , x"FF" , x"E5" , x"C7" , x"A6" , x"A7" , x"EE" , x"B2" , x"FF" , x"DA" , x"B3" , x"E4" , x"C0" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"AA" , x"F6" , x"9F" , x"FD" , x"EE" , x"AF" , x"EB" , x"C1" , x"FF" , x"FD" , x"FF" , x"FD" , x"FF" , x"B3" , x"C0" , x"F2" , x"EB" , x"EC" , x"F1" , x"E2" , x"AF" , x"BC" , x"CC" , x"F0" , x"EA" , x"EA" , x"E9" , x"E8" , x"E8" , x"E7" , x"E7" , x"E7" , x"E6" , x"E4" , x"EA" , x"D5" , x"BB" , x"E9" , x"B0" , x"FF" , x"A1" , x"F6" , x"A5" , x"DE" , x"FE" , x"FD" , x"FF" , x"FD" , x"FE" , x"EC" , x"9B" , x"FC" , x"AA" , x"FF" , x"D4" , x"C2" , x"D6" , x"93" , x"EE" , x"A1" , x"F3" , x"FF" , x"FE" , x"FD" , x"FF" , x"B0" , x"CA" , x"F1" , x"9E" , x"C4" , x"80" , x"79" , x"76" , x"AE" , x"EB" , x"B2" , x"FF" , x"DA" , x"B3" , x"E4" , x"C1" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"AB" , x"F6" , x"A0" , x"FE" , x"EE" , x"AD" , x"EC" , x"C2" , x"FF" , x"FD" , x"FF" , x"FD" , x"FF" , x"A7" , x"ED" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A1" , x"8D" , x"F4" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"FE" , x"FE" , x"FF" , x"FF" , x"FE" , x"FD" , x"FF" , x"E2" , x"C6" , x"E0" , x"BE" , x"FF" , x"A4" , x"FA" , x"A2" , x"FC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A1" , x"F8" , x"AA" , x"FC" , x"E3" , x"B3" , x"E0" , x"96" , x"ED" , x"9F" , x"F1" , x"FF" , x"FE" , x"FD" , x"FF" , x"D5" , x"9C" , x"FA" , x"9F" , x"7F" , x"A5" , x"AA" , x"A2" , x"BE" , x"EA" , x"B1" , x"FF" , x"D9" , x"B1" , x"E4" , x"C1" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"AA" , x"F6" , x"A1" , x"FE" , x"EE" , x"AD" , x"EC" , x"C3" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"A6" , x"F3" , x"D8" , x"D1" , x"D4" , x"CD" , x"F0" , x"B2" , x"9E" , x"F3" , x"D4" , x"D4" , x"D4" , x"D4" , x"D5" , x"D6" , x"D8" , x"D8" , x"D8" , x"DA" , x"D7" , x"E9" , x"D8" , x"C9" , x"D7" , x"C9" , x"FD" , x"A8" , x"F4" , x"AA" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"AA" , x"EC" , x"B1" , x"E9" , x"EC" , x"AB" , x"E4" , x"97" , x"ED" , x"9E" , x"EE" , x"FF" , x"FE" , x"FE" , x"FF" , x"F5" , x"89" , x"F0" , x"C2" , x"A6" , x"F4" , x"F3" , x"F0" , x"F7" , x"ED" , x"AF" , x"FF" , x"D9" , x"B1" , x"E4" , x"C1" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"AA" , x"F6" , x"A0" , x"FE" , x"EC" , x"AE" , x"EB" , x"C3" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"A8" , x"F0" , x"9C" , x"8C" , x"8F" , x"8A" , x"D9" , x"BA" , x"A9" , x"E5" , x"91" , x"8D" , x"8E" , x"8D" , x"8C" , x"8D" , x"8E" , x"8F" , x"90" , x"95" , x"8F" , x"C5" , x"D3" , x"CB" , x"D0" , x"CE" , x"EF" , x"AF" , x"EB" , x"B2" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"B0" , x"DE" , x"BB" , x"DC" , x"F6" , x"A7" , x"E9" , x"99" , x"EC" , x"9C" , x"ED" , x"FF" , x"FE" , x"FF" , x"FE" , x"FF" , x"9F" , x"D7" , x"D3" , x"CA" , x"FF" , x"FC" , x"FD" , x"FF" , x"F3" , x"AE" , x"FF" , x"D8" , x"B2" , x"E4" , x"C0" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"AA" , x"F6" , x"A0" , x"FF" , x"E9" , x"AE" , x"EB" , x"C2" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"A6" , x"F4" , x"96" , x"79" , x"90" , x"8E" , x"E0" , x"BA" , x"A9" , x"EA" , x"97" , x"8A" , x"6B" , x"62" , x"61" , x"62" , x"6C" , x"7D" , x"8E" , x"A2" , x"93" , x"DB" , x"C6" , x"CE" , x"CA" , x"D2" , x"E3" , x"B6" , x"E1" , x"BA" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"B6" , x"D2" , x"C8" , x"CE" , x"FD" , x"A4" , x"EB" , x"9B" , x"EC" , x"9C" , x"EC" , x"FF" , x"FE" , x"FF" , x"FD" , x"FF" , x"C9" , x"C7" , x"D1" , x"D7" , x"D9" , x"C4" , x"C8" , x"CC" , x"C3" , x"B4" , x"FF" , x"D7" , x"B2" , x"E4" , x"BF" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"AA" , x"F6" , x"A0" , x"FF" , x"E7" , x"AD" , x"EA" , x"C2" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"A7" , x"F7" , x"9B" , x"EA" , x"FF" , x"AE" , x"E2" , x"BE" , x"AA" , x"EE" , x"B1" , x"FC" , x"DD" , x"D0" , x"CD" , x"D5" , x"E4" , x"F4" , x"FE" , x"FF" , x"B3" , x"EE" , x"B9" , x"D0" , x"C5" , x"D3" , x"DF" , x"BF" , x"D8" , x"C1" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"C1" , x"C9" , x"D2" , x"C8" , x"FF" , x"9E" , x"EC" , x"9C" , x"EB" , x"9C" , x"EC" , x"FF" , x"FD" , x"FD" , x"FC" , x"FD" , x"DF" , x"C3" , x"D3" , x"D8" , x"AF" , x"89" , x"8E" , x"8E" , x"84" , x"CE" , x"FF" , x"D6" , x"B2" , x"E4" , x"BF" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"AB" , x"F6" , x"A1" , x"FF" , x"E8" , x"AF" , x"EA" , x"C2" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"A8" , x"F8" , x"A5" , x"FF" , x"FF" , x"B2" , x"E1" , x"BE" , x"AA" , x"ED" , x"AB" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"A8" , x"F7" , x"A6" , x"D4" , x"C2" , x"D4" , x"DA" , x"C4" , x"D2" , x"C3" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"C8" , x"C2" , x"D7" , x"C5" , x"FF" , x"9D" , x"ED" , x"9D" , x"EB" , x"9C" , x"EC" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"E6" , x"C3" , x"D2" , x"DC" , x"AF" , x"94" , x"9B" , x"9B" , x"B7" , x"FB" , x"FF" , x"D8" , x"B2" , x"E4" , x"BE" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"AC" , x"F6" , x"9F" , x"FF" , x"E7" , x"AF" , x"EA" , x"C2" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"A8" , x"F8" , x"A3" , x"FE" , x"FF" , x"AF" , x"E1" , x"BD" , x"AA" , x"ED" , x"A7" , x"FE" , x"FD" , x"FE" , x"FD" , x"FC" , x"FD" , x"FC" , x"FE" , x"DC" , x"AE" , x"F3" , x"95" , x"D6" , x"C2" , x"D2" , x"D8" , x"C6" , x"D2" , x"C1" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"CA" , x"C1" , x"D8" , x"C5" , x"FF" , x"9C" , x"ED" , x"9D" , x"EB" , x"9B" , x"EB" , x"FF" , x"F5" , x"BF" , x"B6" , x"B3" , x"92" , x"C7" , x"D3" , x"DF" , x"B4" , x"F7" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"D9" , x"B2" , x"E4" , x"BD" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"AC" , x"F6" , x"9F" , x"FF" , x"E8" , x"B0" , x"EA" , x"C3" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"A9" , x"F8" , x"A5" , x"FF" , x"FF" , x"AC" , x"E1" , x"BE" , x"A9" , x"EE" , x"A7" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"9E" , x"D9" , x"E1" , x"82" , x"D6" , x"C4" , x"CE" , x"DA" , x"C2" , x"D7" , x"BE" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"C8" , x"C4" , x"D4" , x"C7" , x"FF" , x"9C" , x"EC" , x"9C" , x"EB" , x"9A" , x"E9" , x"FF" , x"B2" , x"80" , x"7D" , x"7F" , x"7D" , x"C4" , x"CF" , x"E0" , x"B4" , x"F6" , x"FF" , x"FE" , x"FE" , x"FD" , x"FF" , x"DA" , x"B2" , x"E4" , x"BC" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"AC" , x"F6" , x"9F" , x"FF" , x"E8" , x"B0" , x"EA" , x"C3" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AB" , x"F8" , x"A5" , x"FF" , x"FF" , x"A8" , x"E1" , x"BE" , x"A8" , x"EE" , x"A5" , x"FF" , x"FE" , x"FF" , x"FF" , x"E7" , x"F1" , x"FF" , x"C8" , x"8C" , x"F6" , x"BD" , x"71" , x"D2" , x"C9" , x"C9" , x"DF" , x"BA" , x"DE" , x"B7" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"BF" , x"CE" , x"CD" , x"CB" , x"FA" , x"9F" , x"EB" , x"9C" , x"EB" , x"9A" , x"EA" , x"FF" , x"9C" , x"B4" , x"AD" , x"AE" , x"A6" , x"D5" , x"CC" , x"DE" , x"A7" , x"E0" , x"FF" , x"FE" , x"FF" , x"FE" , x"FF" , x"DB" , x"B2" , x"E4" , x"BC" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"AB" , x"F6" , x"9F" , x"FF" , x"E8" , x"B0" , x"EA" , x"C4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AC" , x"F8" , x"A4" , x"FF" , x"FF" , x"A5" , x"E1" , x"BE" , x"A8" , x"ED" , x"9B" , x"FF" , x"FE" , x"FF" , x"C0" , x"73" , x"81" , x"8B" , x"79" , x"C2" , x"FE" , x"99" , x"9A" , x"CA" , x"D0" , x"C6" , x"E7" , x"AE" , x"E7" , x"B0" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"B4" , x"DB" , x"C1" , x"D4" , x"F1" , x"A3" , x"E8" , x"9A" , x"EC" , x"98" , x"EC" , x"FF" , x"A1" , x"FD" , x"F7" , x"F6" , x"F5" , x"FF" , x"BF" , x"E2" , x"BA" , x"B7" , x"FF" , x"FD" , x"FF" , x"FE" , x"FF" , x"DB" , x"B4" , x"E4" , x"BB" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"AA" , x"F6" , x"9F" , x"FF" , x"E7" , x"B0" , x"EA" , x"C4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AC" , x"F9" , x"A4" , x"FF" , x"FF" , x"A2" , x"E2" , x"BE" , x"A3" , x"F2" , x"8F" , x"EA" , x"FE" , x"FF" , x"8E" , x"91" , x"8A" , x"87" , x"A4" , x"F7" , x"E0" , x"8E" , x"C2" , x"C4" , x"D7" , x"BD" , x"F4" , x"A3" , x"F2" , x"A8" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"AA" , x"E8" , x"B3" , x"E1" , x"E8" , x"A7" , x"E6" , x"99" , x"EC" , x"98" , x"EC" , x"FF" , x"9E" , x"FC" , x"FD" , x"FC" , x"FE" , x"F9" , x"9F" , x"DB" , x"DE" , x"8E" , x"FF" , x"FE" , x"FF" , x"FE" , x"FF" , x"DC" , x"B4" , x"E4" , x"BB" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"A9" , x"F6" , x"9F" , x"FF" , x"E7" , x"B0" , x"EA" , x"C3" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AD" , x"F9" , x"A4" , x"FF" , x"FF" , x"A3" , x"E2" , x"BD" , x"96" , x"FB" , x"B4" , x"B3" , x"FF" , x"FF" , x"95" , x"D5" , x"D2" , x"C6" , x"EC" , x"FF" , x"AC" , x"AA" , x"DB" , x"B9" , x"E1" , x"B0" , x"FE" , x"9A" , x"F8" , x"9F" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"9F" , x"F3" , x"A7" , x"F1" , x"DC" , x"B3" , x"E0" , x"95" , x"ED" , x"9A" , x"EB" , x"FF" , x"9E" , x"F5" , x"C2" , x"BD" , x"C2" , x"B2" , x"81" , x"B6" , x"F6" , x"84" , x"E5" , x"FF" , x"FE" , x"FE" , x"FF" , x"DC" , x"B4" , x"E4" , x"BA" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A8" , x"F6" , x"A0" , x"FF" , x"E7" , x"B0" , x"EA" , x"C4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AD" , x"F9" , x"A5" , x"FF" , x"FF" , x"A4" , x"E2" , x"BC" , x"78" , x"E2" , x"E0" , x"82" , x"FA" , x"FF" , x"95" , x"DE" , x"FF" , x"FC" , x"FF" , x"D5" , x"7B" , x"E8" , x"DF" , x"A9" , x"EA" , x"A4" , x"FF" , x"91" , x"F6" , x"9F" , x"E8" , x"FF" , x"FE" , x"FF" , x"FE" , x"FF" , x"F2" , x"99" , x"F9" , x"9B" , x"FF" , x"CE" , x"C3" , x"D8" , x"92" , x"ED" , x"9A" , x"EB" , x"FF" , x"9C" , x"F0" , x"95" , x"82" , x"88" , x"7E" , x"AE" , x"98" , x"FB" , x"AB" , x"BD" , x"FF" , x"FC" , x"FE" , x"FF" , x"DC" , x"B4" , x"E4" , x"BA" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A5" , x"F6" , x"A0" , x"FF" , x"E7" , x"B0" , x"EA" , x"C4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AD" , x"F9" , x"A5" , x"FF" , x"FF" , x"A8" , x"E3" , x"B8" , x"66" , x"B7" , x"F9" , x"8B" , x"CD" , x"FE" , x"A8" , x"A9" , x"FB" , x"F5" , x"D5" , x"97" , x"9F" , x"FF" , x"DF" , x"A0" , x"F2" , x"99" , x"FF" , x"8D" , x"ED" , x"BD" , x"BF" , x"FF" , x"FD" , x"FF" , x"FD" , x"FE" , x"C8" , x"AD" , x"F5" , x"99" , x"FF" , x"BD" , x"D3" , x"CF" , x"8C" , x"EE" , x"99" , x"EC" , x"FF" , x"9B" , x"F4" , x"9D" , x"AF" , x"AC" , x"D7" , x"FF" , x"96" , x"E8" , x"D5" , x"9B" , x"FF" , x"FE" , x"FE" , x"FF" , x"DC" , x"B3" , x"E4" , x"B9" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A6" , x"F6" , x"9F" , x"FF" , x"E7" , x"B0" , x"E9" , x"C3" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AD" , x"F9" , x"A7" , x"FF" , x"FF" , x"AD" , x"E3" , x"B7" , x"A2" , x"93" , x"F9" , x"BC" , x"97" , x"FF" , x"D4" , x"7A" , x"EF" , x"D2" , x"92" , x"90" , x"EF" , x"FF" , x"ED" , x"98" , x"F7" , x"93" , x"FF" , x"97" , x"D7" , x"E1" , x"8C" , x"FF" , x"FD" , x"FD" , x"FD" , x"FF" , x"90" , x"D4" , x"E4" , x"A1" , x"FF" , x"AC" , x"E4" , x"BC" , x"83" , x"EF" , x"99" , x"EC" , x"FF" , x"9B" , x"F8" , x"A5" , x"FF" , x"FF" , x"FF" , x"FF" , x"B6" , x"C4" , x"F2" , x"8C" , x"F7" , x"FF" , x"FD" , x"FF" , x"DC" , x"B3" , x"E4" , x"B9" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A4" , x"F6" , x"9F" , x"FF" , x"E7" , x"B0" , x"E9" , x"C4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AD" , x"F9" , x"A8" , x"FF" , x"FF" , x"B0" , x"E3" , x"B7" , x"D2" , x"91" , x"E0" , x"E3" , x"7B" , x"F1" , x"FD" , x"7A" , x"CF" , x"EC" , x"8E" , x"E0" , x"FF" , x"FF" , x"FD" , x"94" , x"F6" , x"97" , x"F4" , x"B5" , x"B1" , x"FB" , x"91" , x"BC" , x"FF" , x"FF" , x"FF" , x"CA" , x"86" , x"F5" , x"C0" , x"BC" , x"FF" , x"9B" , x"F2" , x"A4" , x"7B" , x"EF" , x"9B" , x"EC" , x"FF" , x"9E" , x"F8" , x"A3" , x"FD" , x"FE" , x"FC" , x"FF" , x"E0" , x"96" , x"FB" , x"9F" , x"D7" , x"FF" , x"FC" , x"FF" , x"DB" , x"B4" , x"E4" , x"B8" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A4" , x"F6" , x"A1" , x"FF" , x"E6" , x"B0" , x"E9" , x"C5" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AD" , x"F9" , x"A9" , x"FF" , x"FF" , x"B0" , x"E2" , x"B8" , x"DA" , x"BF" , x"B5" , x"FF" , x"96" , x"C0" , x"FF" , x"A9" , x"A2" , x"FF" , x"A5" , x"D4" , x"FE" , x"FD" , x"FF" , x"97" , x"EF" , x"AC" , x"D7" , x"E0" , x"84" , x"FA" , x"C2" , x"73" , x"B9" , x"DF" , x"BA" , x"73" , x"B6" , x"FF" , x"95" , x"E5" , x"FA" , x"90" , x"F9" , x"8E" , x"78" , x"F1" , x"9A" , x"ED" , x"FF" , x"9E" , x"F7" , x"9F" , x"FF" , x"FF" , x"FE" , x"FF" , x"FD" , x"91" , x"ED" , x"CB" , x"B4" , x"FF" , x"FC" , x"FF" , x"DA" , x"B2" , x"E4" , x"B8" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A4" , x"F6" , x"A2" , x"FF" , x"E5" , x"AE" , x"E9" , x"C5" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AC" , x"F9" , x"AA" , x"FF" , x"FF" , x"B1" , x"E2" , x"B7" , x"D5" , x"F3" , x"88" , x"F7" , x"C2" , x"95" , x"FF" , x"E6" , x"7C" , x"EE" , x"D1" , x"A4" , x"FF" , x"FC" , x"FF" , x"9E" , x"DD" , x"CC" , x"B7" , x"FF" , x"79" , x"DA" , x"F4" , x"96" , x"73" , x"70" , x"75" , x"92" , x"ED" , x"E7" , x"8F" , x"FF" , x"D9" , x"9B" , x"F8" , x"96" , x"95" , x"F4" , x"9B" , x"ED" , x"FF" , x"9E" , x"F7" , x"9F" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"AE" , x"CC" , x"EB" , x"9A" , x"FF" , x"FE" , x"FF" , x"D8" , x"B2" , x"E4" , x"B8" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A2" , x"F5" , x"A2" , x"FF" , x"E6" , x"B0" , x"E9" , x"C4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AC" , x"F9" , x"AC" , x"FF" , x"FF" , x"B3" , x"E2" , x"B6" , x"D1" , x"FF" , x"92" , x"DB" , x"E7" , x"7B" , x"F0" , x"FF" , x"92" , x"CB" , x"F1" , x"89" , x"F0" , x"FF" , x"FF" , x"AF" , x"C5" , x"E7" , x"99" , x"FF" , x"A0" , x"A8" , x"FF" , x"DE" , x"9D" , x"8F" , x"9C" , x"D6" , x"FF" , x"B7" , x"A8" , x"FE" , x"B2" , x"BF" , x"ED" , x"A8" , x"A9" , x"F6" , x"9C" , x"ED" , x"FF" , x"9E" , x"F7" , x"A0" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"D6" , x"A0" , x"FB" , x"9A" , x"E9" , x"FF" , x"FF" , x"D7" , x"B3" , x"E4" , x"B9" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A2" , x"F6" , x"A3" , x"FF" , x"E6" , x"B0" , x"E9" , x"C4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AA" , x"F9" , x"AD" , x"FF" , x"FF" , x"B2" , x"E3" , x"B6" , x"D2" , x"FE" , x"BA" , x"AD" , x"FF" , x"96" , x"BD" , x"FE" , x"C5" , x"9D" , x"FF" , x"A9" , x"BE" , x"FF" , x"FF" , x"C6" , x"A5" , x"F6" , x"8B" , x"F6" , x"E3" , x"77" , x"D8" , x"FF" , x"ED" , x"D9" , x"E8" , x"FF" , x"E0" , x"82" , x"DE" , x"FF" , x"8D" , x"DE" , x"D5" , x"B6" , x"AA" , x"F6" , x"9C" , x"ED" , x"FF" , x"9F" , x"F7" , x"9E" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F7" , x"8E" , x"F2" , x"C3" , x"C3" , x"FE" , x"FF" , x"D4" , x"B4" , x"E4" , x"B8" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A2" , x"F6" , x"A4" , x"FF" , x"E4" , x"B0" , x"E9" , x"C4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AC" , x"F9" , x"AD" , x"FF" , x"FF" , x"B3" , x"E2" , x"B6" , x"D4" , x"FF" , x"E8" , x"86" , x"F4" , x"C7" , x"8E" , x"FF" , x"F3" , x"84" , x"EB" , x"D5" , x"89" , x"FF" , x"FF" , x"E1" , x"84" , x"F8" , x"A8" , x"C6" , x"FF" , x"8E" , x"99" , x"E8" , x"FF" , x"FF" , x"FF" , x"EF" , x"A6" , x"90" , x"FF" , x"E5" , x"81" , x"F4" , x"B1" , x"CB" , x"A6" , x"F5" , x"9D" , x"EF" , x"FF" , x"9E" , x"F7" , x"9E" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"A3" , x"D4" , x"E9" , x"A2" , x"FF" , x"FF" , x"D1" , x"B4" , x"E3" , x"B6" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A1" , x"F6" , x"A4" , x"FF" , x"E4" , x"B0" , x"E9" , x"C4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AC" , x"F9" , x"AC" , x"FF" , x"FF" , x"B4" , x"E3" , x"B5" , x"D5" , x"FF" , x"FF" , x"95" , x"D5" , x"EB" , x"7E" , x"E8" , x"FF" , x"A4" , x"C8" , x"F3" , x"81" , x"E2" , x"FF" , x"FC" , x"85" , x"E8" , x"CE" , x"94" , x"FF" , x"DE" , x"6D" , x"9D" , x"D0" , x"E5" , x"D3" , x"A5" , x"72" , x"D7" , x"FF" , x"A8" , x"A7" , x"F9" , x"8E" , x"E5" , x"A1" , x"F4" , x"9E" , x"F1" , x"FF" , x"9E" , x"F7" , x"A0" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"CA" , x"A9" , x"FA" , x"97" , x"ED" , x"FF" , x"CF" , x"B4" , x"E3" , x"B6" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A3" , x"F6" , x"A4" , x"FF" , x"E3" , x"B0" , x"E9" , x"C3" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AB" , x"F9" , x"AA" , x"FF" , x"FF" , x"B6" , x"E3" , x"B5" , x"D6" , x"FF" , x"FF" , x"C5" , x"A6" , x"FF" , x"A1" , x"BC" , x"FE" , x"D0" , x"9A" , x"FD" , x"AC" , x"B4" , x"FF" , x"FF" , x"99" , x"CB" , x"EE" , x"7E" , x"E4" , x"FF" , x"AB" , x"74" , x"8A" , x"95" , x"8C" , x"78" , x"9A" , x"FF" , x"F5" , x"74" , x"D1" , x"EC" , x"8A" , x"FE" , x"98" , x"F4" , x"A0" , x"F2" , x"FF" , x"9B" , x"F7" , x"A1" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F1" , x"8C" , x"F5" , x"BB" , x"C2" , x"FE" , x"CC" , x"B4" , x"E3" , x"B6" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A4" , x"F6" , x"A4" , x"FF" , x"E4" , x"B0" , x"E8" , x"C4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AB" , x"F8" , x"A8" , x"FF" , x"FF" , x"B7" , x"E2" , x"B5" , x"D7" , x"FF" , x"FF" , x"F3" , x"8A" , x"F1" , x"CD" , x"91" , x"FF" , x"F8" , x"8A" , x"EA" , x"D7" , x"8C" , x"FE" , x"FF" , x"C0" , x"A0" , x"FF" , x"AA" , x"A0" , x"FF" , x"FE" , x"A5" , x"67" , x"70" , x"62" , x"8D" , x"F7" , x"FF" , x"B6" , x"88" , x"F5" , x"CB" , x"A0" , x"FF" , x"92" , x"F4" , x"9E" , x"F1" , x"FF" , x"9A" , x"F7" , x"A2" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"9F" , x"DD" , x"E2" , x"98" , x"FF" , x"CC" , x"B4" , x"E3" , x"B7" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A2" , x"F6" , x"A2" , x"FF" , x"E4" , x"B0" , x"E8" , x"C4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AB" , x"F9" , x"A7" , x"FF" , x"FF" , x"B8" , x"E3" , x"B5" , x"D7" , x"FF" , x"FC" , x"FF" , x"A4" , x"D1" , x"F0" , x"7F" , x"E9" , x"FF" , x"AD" , x"C2" , x"F6" , x"84" , x"DA" , x"FE" , x"E9" , x"7E" , x"EE" , x"D8" , x"75" , x"DB" , x"FF" , x"FF" , x"DA" , x"B7" , x"CD" , x"FF" , x"FF" , x"F1" , x"70" , x"B4" , x"FF" , x"9D" , x"C7" , x"FF" , x"92" , x"F3" , x"9D" , x"F0" , x"FF" , x"9A" , x"F7" , x"A5" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FE" , x"C6" , x"B3" , x"F8" , x"8C" , x"F6" , x"D2" , x"B5" , x"E3" , x"B7" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A4" , x"F6" , x"A1" , x"FE" , x"E4" , x"B1" , x"E7" , x"C4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AC" , x"F9" , x"A6" , x"FE" , x"FD" , x"B9" , x"E2" , x"B5" , x"D7" , x"FF" , x"FB" , x"FE" , x"CF" , x"A2" , x"FF" , x"A5" , x"B7" , x"FE" , x"DF" , x"92" , x"FD" , x"B2" , x"A3" , x"FF" , x"FF" , x"8B" , x"C6" , x"FF" , x"A0" , x"85" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"9B" , x"87" , x"E8" , x"E6" , x"7B" , x"F0" , x"FF" , x"94" , x"F3" , x"9B" , x"EC" , x"FE" , x"99" , x"F7" , x"A5" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"ED" , x"8F" , x"F9" , x"B5" , x"CC" , x"D8" , x"B6" , x"E3" , x"B6" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A4" , x"F6" , x"9F" , x"FF" , x"E5" , x"B1" , x"E7" , x"C5" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AC" , x"F9" , x"A6" , x"FF" , x"FF" , x"BB" , x"E3" , x"B5" , x"D6" , x"FF" , x"FD" , x"FF" , x"F6" , x"8B" , x"ED" , x"D2" , x"86" , x"FF" , x"FE" , x"95" , x"E6" , x"DC" , x"7B" , x"F3" , x"FF" , x"BB" , x"93" , x"FA" , x"D7" , x"83" , x"97" , x"E7" , x"FF" , x"FF" , x"FF" , x"ED" , x"A3" , x"70" , x"B9" , x"FF" , x"B6" , x"90" , x"FF" , x"FF" , x"97" , x"F3" , x"98" , x"ED" , x"FF" , x"95" , x"F7" , x"A5" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"9D" , x"E3" , x"DC" , x"9D" , x"D0" , x"B7" , x"E3" , x"B4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A4" , x"F2" , x"97" , x"F4" , x"DD" , x"B0" , x"E5" , x"C9" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AB" , x"F6" , x"95" , x"B2" , x"BD" , x"8D" , x"E1" , x"B5" , x"D7" , x"FF" , x"FD" , x"FE" , x"FF" , x"A7" , x"CA" , x"F4" , x"80" , x"C6" , x"FF" , x"99" , x"C2" , x"F8" , x"8B" , x"C7" , x"FF" , x"F0" , x"78" , x"CD" , x"FF" , x"B3" , x"7C" , x"68" , x"7A" , x"80" , x"77" , x"64" , x"71" , x"9A" , x"F2" , x"EB" , x"84" , x"C9" , x"FF" , x"FF" , x"9A" , x"F2" , x"93" , x"D2" , x"E0" , x"88" , x"F6" , x"A5" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FE" , x"BF" , x"BC" , x"F5" , x"89" , x"95" , x"B6" , x"E3" , x"B4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"A6" , x"F0" , x"99" , x"8C" , x"87" , x"BA" , x"E1" , x"CD" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"AD" , x"F3" , x"97" , x"75" , x"75" , x"7E" , x"DD" , x"B4" , x"DA" , x"FF" , x"FE" , x"FD" , x"FF" , x"D3" , x"98" , x"FD" , x"AA" , x"70" , x"8C" , x"80" , x"A4" , x"FA" , x"B8" , x"A6" , x"FF" , x"FF" , x"A5" , x"98" , x"F1" , x"F3" , x"AC" , x"83" , x"78" , x"77" , x"77" , x"7F" , x"98" , x"E0" , x"FF" , x"B6" , x"81" , x"FB" , x"FF" , x"FF" , x"9D" , x"EF" , x"9E" , x"78" , x"76" , x"92" , x"F2" , x"A5" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"E5" , x"93" , x"FA" , x"A5" , x"6B" , x"BD" , x"E3" , x"B4" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"A6" , x"F1" , x"A9" , x"8A" , x"85" , x"CC" , x"D7" , x"D3" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"AE" , x"F1" , x"A1" , x"95" , x"99" , x"91" , x"DE" , x"B6" , x"E0" , x"FF" , x"FE" , x"FF" , x"FF" , x"F8" , x"88" , x"EB" , x"D3" , x"86" , x"8E" , x"91" , x"8F" , x"DC" , x"E2" , x"9F" , x"FF" , x"FE" , x"EB" , x"75" , x"BC" , x"FD" , x"F0" , x"BB" , x"9A" , x"97" , x"99" , x"AD" , x"E3" , x"FF" , x"D5" , x"7F" , x"D1" , x"FF" , x"FD" , x"FF" , x"A0" , x"EE" , x"A6" , x"89" , x"88" , x"9B" , x"F1" , x"A8" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"95" , x"EB" , x"D0" , x"7E" , x"BE" , x"E3" , x"B9" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"A8" , x"E9" , x"E4" , x"D4" , x"CF" , x"F0" , x"BF" , x"DD" , x"FF" , x"FE" , x"FF" , x"FE" , x"FF" , x"AD" , x"F4" , x"E6" , x"E1" , x"E2" , x"DE" , x"F9" , x"B1" , x"E8" , x"FF" , x"FE" , x"FF" , x"FE" , x"FF" , x"A4" , x"C2" , x"F9" , x"CF" , x"D5" , x"D4" , x"D0" , x"E7" , x"EA" , x"A7" , x"FF" , x"FC" , x"FF" , x"B3" , x"87" , x"D2" , x"FF" , x"FC" , x"E9" , x"E1" , x"E5" , x"F5" , x"FF" , x"E9" , x"9A" , x"99" , x"FF" , x"FE" , x"FE" , x"FF" , x"A4" , x"ED" , x"E0" , x"D3" , x"D4" , x"DB" , x"F4" , x"AB" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"B4" , x"C7" , x"F7" , x"CC" , x"EC" , x"D9" , x"BC" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"AF" , x"D3" , x"FF" , x"FE" , x"FD" , x"FF" , x"A8" , x"EE" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"AD" , x"E7" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"A3" , x"F7" , x"FF" , x"FE" , x"FF" , x"FD" , x"FF" , x"D6" , x"91" , x"F7" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"E9" , x"AB" , x"FF" , x"FC" , x"FE" , x"FA" , x"88" , x"93" , x"D1" , x"FB" , x"FF" , x"FF" , x"FF" , x"FE" , x"E1" , x"A2" , x"82" , x"EE" , x"FE" , x"FE" , x"FD" , x"FF" , x"AB" , x"DB" , x"FF" , x"FD" , x"FF" , x"FF" , x"E6" , x"AA" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"DC" , x"9B" , x"FC" , x"FF" , x"FF" , x"C0" , x"C7" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"CA" , x"A6" , x"EC" , x"E8" , x"EE" , x"DD" , x"9F" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"C0" , x"B5" , x"E6" , x"DD" , x"DE" , x"E5" , x"D2" , x"9D" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FB" , x"8D" , x"DB" , x"F2" , x"EB" , x"EA" , x"EA" , x"F1" , x"DF" , x"B6" , x"FF" , x"FD" , x"FE" , x"FF" , x"E8" , x"7A" , x"8D" , x"B2" , x"D5" , x"DF" , x"DB" , x"C1" , x"96" , x"79" , x"D4" , x"FF" , x"FE" , x"FF" , x"FD" , x"FF" , x"C2" , x"AC" , x"EC" , x"E8" , x"E8" , x"EC" , x"B5" , x"BD" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FB" , x"91" , x"E0" , x"EE" , x"E3" , x"93" , x"E5" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F0" , x"7E" , x"9E" , x"A0" , x"A0" , x"98" , x"C5" , x"FF" , x"FE" , x"FF" , x"FF" , x"FE" , x"FF" , x"EA" , x"81" , x"95" , x"92" , x"93" , x"94" , x"8D" , x"C9" , x"FF" , x"FD" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"B6" , x"9C" , x"A4" , x"9F" , x"9F" , x"9F" , x"A2" , x"9A" , x"CB" , x"FF" , x"FD" , x"FF" , x"FE" , x"FF" , x"DC" , x"7E" , x"7F" , x"8D" , x"93" , x"91" , x"86" , x"7D" , x"CD" , x"FF" , x"FD" , x"FF" , x"FF" , x"FD" , x"FF" , x"E9" , x"7A" , x"9F" , x"A0" , x"A0" , x"9D" , x"83" , x"EA" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FF" , x"B9" , x"9A" , x"A2" , x"9C" , x"99" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"C0" , x"76" , x"7A" , x"7D" , x"A4" , x"FA" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"C7" , x"89" , x"7C" , x"7B" , x"87" , x"B5" , x"FE" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FD" , x"FE" , x"EE" , x"7C" , x"80" , x"7B" , x"7C" , x"7B" , x"7E" , x"83" , x"F0" , x"FF" , x"FE" , x"FF" , x"FF" , x"FE" , x"FF" , x"F0" , x"A4" , x"7A" , x"78" , x"81" , x"A8" , x"E9" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"A8" , x"79" , x"7D" , x"7D" , x"76" , x"C1" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FE" , x"F1" , x"86" , x"80" , x"7B" , x"E1" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"D7" , x"C6" , x"DB" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"F8" , x"ED" , x"EE" , x"F6" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"D6" , x"9A" , x"A2" , x"AF" , x"B4" , x"B9" , x"E7" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"F3" , x"E8" , x"F3" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FF" , x"BF" , x"A3" , x"AB" , x"D0" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"E8" , x"AB" , x"DA" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FE" , x"FE" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"FD" , x"FD" , x"FD" , x"FD" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FD" , x"FD" , x"FD" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FE" , x"FD" , x"FE" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ),
( x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" , x"FF" ) 
);

END PACKAGE texturas;

-------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------------

PACKAGE BODY texturas IS

END texturas;